
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"a6",x"c4",x"87",x"c7"),
     1 => (x"c5",x"78",x"c0",x"48"),
     2 => (x"48",x"a6",x"c4",x"87"),
     3 => (x"66",x"c4",x"78",x"c1"),
     4 => (x"ee",x"49",x"73",x"1e"),
     5 => (x"86",x"c8",x"87",x"df"),
     6 => (x"ef",x"49",x"e0",x"c0"),
     7 => (x"a5",x"c4",x"87",x"ef"),
     8 => (x"f0",x"49",x"6a",x"4a"),
     9 => (x"c6",x"f1",x"87",x"f0"),
    10 => (x"c1",x"85",x"cb",x"87"),
    11 => (x"ab",x"b7",x"c8",x"83"),
    12 => (x"87",x"c7",x"ff",x"04"),
    13 => (x"26",x"4d",x"26",x"26"),
    14 => (x"26",x"4b",x"26",x"4c"),
    15 => (x"4a",x"71",x"1e",x"4f"),
    16 => (x"5a",x"f2",x"f0",x"c2"),
    17 => (x"48",x"f2",x"f0",x"c2"),
    18 => (x"fe",x"49",x"78",x"c7"),
    19 => (x"4f",x"26",x"87",x"dd"),
    20 => (x"71",x"1e",x"73",x"1e"),
    21 => (x"aa",x"b7",x"c0",x"4a"),
    22 => (x"c2",x"87",x"d3",x"03"),
    23 => (x"05",x"bf",x"dd",x"d1"),
    24 => (x"4b",x"c1",x"87",x"c4"),
    25 => (x"4b",x"c0",x"87",x"c2"),
    26 => (x"5b",x"e1",x"d1",x"c2"),
    27 => (x"d1",x"c2",x"87",x"c4"),
    28 => (x"d1",x"c2",x"5a",x"e1"),
    29 => (x"c1",x"4a",x"bf",x"dd"),
    30 => (x"a2",x"c0",x"c1",x"9a"),
    31 => (x"87",x"e8",x"ec",x"49"),
    32 => (x"bf",x"c5",x"d1",x"c2"),
    33 => (x"dd",x"d1",x"c2",x"49"),
    34 => (x"48",x"fc",x"b1",x"bf"),
    35 => (x"e8",x"fe",x"78",x"71"),
    36 => (x"4a",x"71",x"1e",x"87"),
    37 => (x"72",x"1e",x"66",x"c4"),
    38 => (x"87",x"ee",x"e9",x"49"),
    39 => (x"1e",x"4f",x"26",x"26"),
    40 => (x"bf",x"dd",x"d1",x"c2"),
    41 => (x"87",x"c8",x"e6",x"49"),
    42 => (x"48",x"e6",x"f0",x"c2"),
    43 => (x"c2",x"78",x"bf",x"e8"),
    44 => (x"ec",x"48",x"e2",x"f0"),
    45 => (x"f0",x"c2",x"78",x"bf"),
    46 => (x"49",x"4a",x"bf",x"e6"),
    47 => (x"c8",x"99",x"ff",x"c3"),
    48 => (x"48",x"72",x"2a",x"b7"),
    49 => (x"f0",x"c2",x"b0",x"71"),
    50 => (x"4f",x"26",x"58",x"ee"),
    51 => (x"5c",x"5b",x"5e",x"0e"),
    52 => (x"4b",x"71",x"0e",x"5d"),
    53 => (x"c2",x"87",x"c8",x"ff"),
    54 => (x"c0",x"48",x"e1",x"f0"),
    55 => (x"e5",x"49",x"73",x"50"),
    56 => (x"49",x"70",x"87",x"ee"),
    57 => (x"cb",x"9c",x"c2",x"4c"),
    58 => (x"f8",x"cd",x"49",x"ee"),
    59 => (x"4d",x"49",x"70",x"87"),
    60 => (x"97",x"e1",x"f0",x"c2"),
    61 => (x"e2",x"c1",x"05",x"bf"),
    62 => (x"49",x"66",x"d0",x"87"),
    63 => (x"bf",x"ea",x"f0",x"c2"),
    64 => (x"87",x"d6",x"05",x"99"),
    65 => (x"c2",x"49",x"66",x"d4"),
    66 => (x"99",x"bf",x"e2",x"f0"),
    67 => (x"73",x"87",x"cb",x"05"),
    68 => (x"87",x"fc",x"e4",x"49"),
    69 => (x"c1",x"02",x"98",x"70"),
    70 => (x"4c",x"c1",x"87",x"c1"),
    71 => (x"75",x"87",x"c0",x"fe"),
    72 => (x"87",x"cd",x"cd",x"49"),
    73 => (x"c6",x"02",x"98",x"70"),
    74 => (x"e1",x"f0",x"c2",x"87"),
    75 => (x"c2",x"50",x"c1",x"48"),
    76 => (x"bf",x"97",x"e1",x"f0"),
    77 => (x"87",x"e3",x"c0",x"05"),
    78 => (x"bf",x"ea",x"f0",x"c2"),
    79 => (x"99",x"66",x"d0",x"49"),
    80 => (x"87",x"d6",x"ff",x"05"),
    81 => (x"bf",x"e2",x"f0",x"c2"),
    82 => (x"99",x"66",x"d4",x"49"),
    83 => (x"87",x"ca",x"ff",x"05"),
    84 => (x"fb",x"e3",x"49",x"73"),
    85 => (x"05",x"98",x"70",x"87"),
    86 => (x"74",x"87",x"ff",x"fe"),
    87 => (x"87",x"d5",x"fb",x"48"),
    88 => (x"5c",x"5b",x"5e",x"0e"),
    89 => (x"86",x"f8",x"0e",x"5d"),
    90 => (x"ec",x"4c",x"4d",x"c0"),
    91 => (x"a6",x"c4",x"7e",x"bf"),
    92 => (x"ee",x"f0",x"c2",x"48"),
    93 => (x"1e",x"c0",x"78",x"bf"),
    94 => (x"49",x"f7",x"c1",x"1e"),
    95 => (x"c8",x"87",x"cd",x"fd"),
    96 => (x"02",x"98",x"70",x"86"),
    97 => (x"c2",x"87",x"f3",x"c0"),
    98 => (x"05",x"bf",x"c5",x"d1"),
    99 => (x"7e",x"c1",x"87",x"c4"),
   100 => (x"7e",x"c0",x"87",x"c2"),
   101 => (x"48",x"c5",x"d1",x"c2"),
   102 => (x"fc",x"ca",x"78",x"6e"),
   103 => (x"02",x"66",x"c4",x"1e"),
   104 => (x"a6",x"c4",x"87",x"c9"),
   105 => (x"dc",x"cf",x"c2",x"48"),
   106 => (x"c4",x"87",x"c7",x"78"),
   107 => (x"cf",x"c2",x"48",x"a6"),
   108 => (x"66",x"c4",x"78",x"e7"),
   109 => (x"87",x"fb",x"c8",x"49"),
   110 => (x"1e",x"c1",x"86",x"c4"),
   111 => (x"49",x"c7",x"1e",x"c0"),
   112 => (x"c8",x"87",x"c9",x"fc"),
   113 => (x"02",x"98",x"70",x"86"),
   114 => (x"49",x"ff",x"87",x"cd"),
   115 => (x"c1",x"87",x"c1",x"fa"),
   116 => (x"fb",x"e1",x"49",x"da"),
   117 => (x"c2",x"4d",x"c1",x"87"),
   118 => (x"bf",x"97",x"e1",x"f0"),
   119 => (x"d6",x"87",x"c3",x"02"),
   120 => (x"f0",x"c2",x"87",x"ef"),
   121 => (x"c2",x"4b",x"bf",x"e6"),
   122 => (x"05",x"bf",x"dd",x"d1"),
   123 => (x"c2",x"87",x"e1",x"c1"),
   124 => (x"02",x"bf",x"c5",x"d1"),
   125 => (x"c4",x"87",x"f0",x"c0"),
   126 => (x"c0",x"c8",x"48",x"a6"),
   127 => (x"d1",x"c2",x"78",x"c0"),
   128 => (x"97",x"6e",x"7e",x"c9"),
   129 => (x"48",x"6e",x"49",x"bf"),
   130 => (x"7e",x"70",x"80",x"c1"),
   131 => (x"87",x"c0",x"e1",x"71"),
   132 => (x"c3",x"02",x"98",x"70"),
   133 => (x"b3",x"66",x"c4",x"87"),
   134 => (x"c1",x"48",x"66",x"c4"),
   135 => (x"a6",x"c8",x"28",x"b7"),
   136 => (x"05",x"98",x"70",x"58"),
   137 => (x"c3",x"87",x"db",x"ff"),
   138 => (x"e3",x"e0",x"49",x"fd"),
   139 => (x"49",x"fa",x"c3",x"87"),
   140 => (x"73",x"87",x"dd",x"e0"),
   141 => (x"99",x"ff",x"c3",x"49"),
   142 => (x"49",x"c0",x"1e",x"71"),
   143 => (x"73",x"87",x"d2",x"f9"),
   144 => (x"29",x"b7",x"c8",x"49"),
   145 => (x"49",x"c1",x"1e",x"71"),
   146 => (x"c8",x"87",x"c6",x"f9"),
   147 => (x"87",x"c7",x"c6",x"86"),
   148 => (x"bf",x"ea",x"f0",x"c2"),
   149 => (x"df",x"02",x"9b",x"4b"),
   150 => (x"d9",x"d1",x"c2",x"87"),
   151 => (x"d0",x"c8",x"49",x"bf"),
   152 => (x"05",x"98",x"70",x"87"),
   153 => (x"c0",x"87",x"c4",x"c0"),
   154 => (x"c2",x"87",x"d3",x"4b"),
   155 => (x"f4",x"c7",x"49",x"e0"),
   156 => (x"dd",x"d1",x"c2",x"87"),
   157 => (x"87",x"c6",x"c0",x"58"),
   158 => (x"48",x"d9",x"d1",x"c2"),
   159 => (x"49",x"73",x"78",x"c0"),
   160 => (x"c0",x"05",x"99",x"c2"),
   161 => (x"eb",x"c3",x"87",x"cf"),
   162 => (x"c3",x"df",x"ff",x"49"),
   163 => (x"c2",x"49",x"70",x"87"),
   164 => (x"c2",x"c0",x"02",x"99"),
   165 => (x"73",x"4c",x"fb",x"87"),
   166 => (x"05",x"99",x"c1",x"49"),
   167 => (x"c3",x"87",x"cf",x"c0"),
   168 => (x"de",x"ff",x"49",x"f4"),
   169 => (x"49",x"70",x"87",x"ea"),
   170 => (x"c0",x"02",x"99",x"c2"),
   171 => (x"4c",x"fa",x"87",x"c2"),
   172 => (x"99",x"c8",x"49",x"73"),
   173 => (x"87",x"cf",x"c0",x"05"),
   174 => (x"ff",x"49",x"f5",x"c3"),
   175 => (x"70",x"87",x"d1",x"de"),
   176 => (x"02",x"99",x"c2",x"49"),
   177 => (x"c2",x"87",x"d6",x"c0"),
   178 => (x"02",x"bf",x"f2",x"f0"),
   179 => (x"48",x"87",x"ca",x"c0"),
   180 => (x"f0",x"c2",x"88",x"c1"),
   181 => (x"c2",x"c0",x"58",x"f6"),
   182 => (x"c1",x"4c",x"ff",x"87"),
   183 => (x"c4",x"49",x"73",x"4d"),
   184 => (x"cf",x"c0",x"05",x"99"),
   185 => (x"49",x"f2",x"c3",x"87"),
   186 => (x"87",x"e4",x"dd",x"ff"),
   187 => (x"99",x"c2",x"49",x"70"),
   188 => (x"87",x"dc",x"c0",x"02"),
   189 => (x"bf",x"f2",x"f0",x"c2"),
   190 => (x"b7",x"c7",x"48",x"7e"),
   191 => (x"cb",x"c0",x"03",x"a8"),
   192 => (x"c1",x"48",x"6e",x"87"),
   193 => (x"f6",x"f0",x"c2",x"80"),
   194 => (x"87",x"c2",x"c0",x"58"),
   195 => (x"4d",x"c1",x"4c",x"fe"),
   196 => (x"ff",x"49",x"fd",x"c3"),
   197 => (x"70",x"87",x"f9",x"dc"),
   198 => (x"02",x"99",x"c2",x"49"),
   199 => (x"c2",x"87",x"d5",x"c0"),
   200 => (x"02",x"bf",x"f2",x"f0"),
   201 => (x"c2",x"87",x"c9",x"c0"),
   202 => (x"c0",x"48",x"f2",x"f0"),
   203 => (x"87",x"c2",x"c0",x"78"),
   204 => (x"4d",x"c1",x"4c",x"fd"),
   205 => (x"ff",x"49",x"fa",x"c3"),
   206 => (x"70",x"87",x"d5",x"dc"),
   207 => (x"02",x"99",x"c2",x"49"),
   208 => (x"c2",x"87",x"d9",x"c0"),
   209 => (x"48",x"bf",x"f2",x"f0"),
   210 => (x"03",x"a8",x"b7",x"c7"),
   211 => (x"c2",x"87",x"c9",x"c0"),
   212 => (x"c7",x"48",x"f2",x"f0"),
   213 => (x"87",x"c2",x"c0",x"78"),
   214 => (x"4d",x"c1",x"4c",x"fc"),
   215 => (x"03",x"ac",x"b7",x"c0"),
   216 => (x"c4",x"87",x"d5",x"c0"),
   217 => (x"d8",x"c1",x"48",x"66"),
   218 => (x"6e",x"7e",x"70",x"80"),
   219 => (x"c7",x"c0",x"02",x"bf"),
   220 => (x"4b",x"bf",x"6e",x"87"),
   221 => (x"0f",x"73",x"49",x"74"),
   222 => (x"f0",x"c3",x"1e",x"c0"),
   223 => (x"49",x"da",x"c1",x"1e"),
   224 => (x"c8",x"87",x"c9",x"f5"),
   225 => (x"02",x"98",x"70",x"86"),
   226 => (x"c2",x"87",x"d9",x"c0"),
   227 => (x"7e",x"bf",x"f2",x"f0"),
   228 => (x"91",x"cb",x"49",x"6e"),
   229 => (x"71",x"4a",x"66",x"c4"),
   230 => (x"c0",x"02",x"6a",x"82"),
   231 => (x"4b",x"6a",x"87",x"c6"),
   232 => (x"0f",x"73",x"49",x"6e"),
   233 => (x"c0",x"02",x"9d",x"75"),
   234 => (x"f0",x"c2",x"87",x"c8"),
   235 => (x"f0",x"49",x"bf",x"f2"),
   236 => (x"d1",x"c2",x"87",x"f9"),
   237 => (x"c0",x"02",x"bf",x"e1"),
   238 => (x"c2",x"49",x"87",x"dd"),
   239 => (x"98",x"70",x"87",x"f3"),
   240 => (x"87",x"d3",x"c0",x"02"),
   241 => (x"bf",x"f2",x"f0",x"c2"),
   242 => (x"87",x"df",x"f0",x"49"),
   243 => (x"ff",x"f1",x"49",x"c0"),
   244 => (x"e1",x"d1",x"c2",x"87"),
   245 => (x"f8",x"78",x"c0",x"48"),
   246 => (x"87",x"d9",x"f1",x"8e"),
   247 => (x"6b",x"79",x"6f",x"4a"),
   248 => (x"20",x"73",x"79",x"65"),
   249 => (x"4a",x"00",x"6e",x"6f"),
   250 => (x"65",x"6b",x"79",x"6f"),
   251 => (x"6f",x"20",x"73",x"79"),
   252 => (x"0e",x"00",x"66",x"66"),
   253 => (x"5d",x"5c",x"5b",x"5e"),
   254 => (x"4c",x"71",x"1e",x"0e"),
   255 => (x"bf",x"ee",x"f0",x"c2"),
   256 => (x"a1",x"cd",x"c1",x"49"),
   257 => (x"81",x"d1",x"c1",x"4d"),
   258 => (x"9c",x"74",x"7e",x"69"),
   259 => (x"c4",x"87",x"cf",x"02"),
   260 => (x"7b",x"74",x"4b",x"a5"),
   261 => (x"bf",x"ee",x"f0",x"c2"),
   262 => (x"87",x"e1",x"f0",x"49"),
   263 => (x"9c",x"74",x"7b",x"6e"),
   264 => (x"c0",x"87",x"c4",x"05"),
   265 => (x"c1",x"87",x"c2",x"4b"),
   266 => (x"f0",x"49",x"73",x"4b"),
   267 => (x"66",x"d4",x"87",x"e2"),
   268 => (x"49",x"87",x"c8",x"02"),
   269 => (x"70",x"87",x"ee",x"c0"),
   270 => (x"c0",x"87",x"c2",x"4a"),
   271 => (x"e5",x"d1",x"c2",x"4a"),
   272 => (x"f0",x"ef",x"26",x"5a"),
   273 => (x"00",x"00",x"00",x"87"),
   274 => (x"11",x"12",x"58",x"00"),
   275 => (x"1c",x"1b",x"1d",x"14"),
   276 => (x"91",x"59",x"5a",x"23"),
   277 => (x"eb",x"f2",x"f5",x"94"),
   278 => (x"00",x"00",x"00",x"f4"),
   279 => (x"00",x"00",x"00",x"00"),
   280 => (x"00",x"00",x"00",x"00"),
   281 => (x"4a",x"71",x"1e",x"00"),
   282 => (x"49",x"bf",x"c8",x"ff"),
   283 => (x"26",x"48",x"a1",x"72"),
   284 => (x"c8",x"ff",x"1e",x"4f"),
   285 => (x"c0",x"fe",x"89",x"bf"),
   286 => (x"c0",x"c0",x"c0",x"c0"),
   287 => (x"87",x"c4",x"01",x"a9"),
   288 => (x"87",x"c2",x"4a",x"c0"),
   289 => (x"48",x"72",x"4a",x"c1"),
   290 => (x"5e",x"0e",x"4f",x"26"),
   291 => (x"0e",x"5d",x"5c",x"5b"),
   292 => (x"d4",x"ff",x"4b",x"71"),
   293 => (x"48",x"66",x"d0",x"4c"),
   294 => (x"49",x"d6",x"78",x"c0"),
   295 => (x"87",x"f0",x"d8",x"ff"),
   296 => (x"6c",x"7c",x"ff",x"c3"),
   297 => (x"99",x"ff",x"c3",x"49"),
   298 => (x"c3",x"49",x"4d",x"71"),
   299 => (x"e0",x"c1",x"99",x"f0"),
   300 => (x"87",x"cb",x"05",x"a9"),
   301 => (x"6c",x"7c",x"ff",x"c3"),
   302 => (x"d0",x"98",x"c3",x"48"),
   303 => (x"c3",x"78",x"08",x"66"),
   304 => (x"4a",x"6c",x"7c",x"ff"),
   305 => (x"c3",x"31",x"c8",x"49"),
   306 => (x"4a",x"6c",x"7c",x"ff"),
   307 => (x"49",x"72",x"b2",x"71"),
   308 => (x"ff",x"c3",x"31",x"c8"),
   309 => (x"71",x"4a",x"6c",x"7c"),
   310 => (x"c8",x"49",x"72",x"b2"),
   311 => (x"7c",x"ff",x"c3",x"31"),
   312 => (x"b2",x"71",x"4a",x"6c"),
   313 => (x"c0",x"48",x"d0",x"ff"),
   314 => (x"9b",x"73",x"78",x"e0"),
   315 => (x"72",x"87",x"c2",x"02"),
   316 => (x"26",x"48",x"75",x"7b"),
   317 => (x"26",x"4c",x"26",x"4d"),
   318 => (x"1e",x"4f",x"26",x"4b"),
   319 => (x"5e",x"0e",x"4f",x"26"),
   320 => (x"f8",x"0e",x"5c",x"5b"),
   321 => (x"c8",x"1e",x"76",x"86"),
   322 => (x"fd",x"fd",x"49",x"a6"),
   323 => (x"70",x"86",x"c4",x"87"),
   324 => (x"c2",x"48",x"6e",x"4b"),
   325 => (x"c6",x"c3",x"03",x"a8"),
   326 => (x"c3",x"4a",x"73",x"87"),
   327 => (x"d0",x"c1",x"9a",x"f0"),
   328 => (x"87",x"c7",x"02",x"aa"),
   329 => (x"05",x"aa",x"e0",x"c1"),
   330 => (x"73",x"87",x"f4",x"c2"),
   331 => (x"02",x"99",x"c8",x"49"),
   332 => (x"c6",x"ff",x"87",x"c3"),
   333 => (x"c3",x"4c",x"73",x"87"),
   334 => (x"05",x"ac",x"c2",x"9c"),
   335 => (x"c4",x"87",x"cd",x"c1"),
   336 => (x"31",x"c9",x"49",x"66"),
   337 => (x"66",x"c4",x"1e",x"71"),
   338 => (x"c2",x"92",x"d4",x"4a"),
   339 => (x"72",x"49",x"f6",x"f0"),
   340 => (x"da",x"d1",x"fe",x"81"),
   341 => (x"49",x"66",x"c4",x"87"),
   342 => (x"49",x"e3",x"c0",x"1e"),
   343 => (x"87",x"d5",x"d6",x"ff"),
   344 => (x"d5",x"ff",x"49",x"d8"),
   345 => (x"c0",x"c8",x"87",x"ea"),
   346 => (x"e6",x"df",x"c2",x"1e"),
   347 => (x"ea",x"ed",x"fd",x"49"),
   348 => (x"48",x"d0",x"ff",x"87"),
   349 => (x"c2",x"78",x"e0",x"c0"),
   350 => (x"d0",x"1e",x"e6",x"df"),
   351 => (x"92",x"d4",x"4a",x"66"),
   352 => (x"49",x"f6",x"f0",x"c2"),
   353 => (x"cf",x"fe",x"81",x"72"),
   354 => (x"86",x"d0",x"87",x"e2"),
   355 => (x"c1",x"05",x"ac",x"c1"),
   356 => (x"66",x"c4",x"87",x"cd"),
   357 => (x"71",x"31",x"c9",x"49"),
   358 => (x"4a",x"66",x"c4",x"1e"),
   359 => (x"f0",x"c2",x"92",x"d4"),
   360 => (x"81",x"72",x"49",x"f6"),
   361 => (x"87",x"c7",x"d0",x"fe"),
   362 => (x"1e",x"e6",x"df",x"c2"),
   363 => (x"d4",x"4a",x"66",x"c8"),
   364 => (x"f6",x"f0",x"c2",x"92"),
   365 => (x"fe",x"81",x"72",x"49"),
   366 => (x"c8",x"87",x"ee",x"cd"),
   367 => (x"c0",x"1e",x"49",x"66"),
   368 => (x"d4",x"ff",x"49",x"e3"),
   369 => (x"49",x"d7",x"87",x"ef"),
   370 => (x"87",x"c4",x"d4",x"ff"),
   371 => (x"c2",x"1e",x"c0",x"c8"),
   372 => (x"fd",x"49",x"e6",x"df"),
   373 => (x"d0",x"87",x"ee",x"eb"),
   374 => (x"48",x"d0",x"ff",x"86"),
   375 => (x"f8",x"78",x"e0",x"c0"),
   376 => (x"87",x"d1",x"fc",x"8e"),
   377 => (x"5c",x"5b",x"5e",x"0e"),
   378 => (x"71",x"1e",x"0e",x"5d"),
   379 => (x"4c",x"d4",x"ff",x"4d"),
   380 => (x"48",x"7e",x"66",x"d4"),
   381 => (x"06",x"a8",x"b7",x"c3"),
   382 => (x"48",x"c0",x"87",x"c5"),
   383 => (x"75",x"87",x"e2",x"c1"),
   384 => (x"fb",x"dd",x"fe",x"49"),
   385 => (x"c4",x"1e",x"75",x"87"),
   386 => (x"93",x"d4",x"4b",x"66"),
   387 => (x"83",x"f6",x"f0",x"c2"),
   388 => (x"c8",x"fe",x"49",x"73"),
   389 => (x"83",x"c8",x"87",x"f7"),
   390 => (x"d0",x"ff",x"4b",x"6b"),
   391 => (x"78",x"e1",x"c8",x"48"),
   392 => (x"49",x"73",x"7c",x"dd"),
   393 => (x"71",x"99",x"ff",x"c3"),
   394 => (x"c8",x"49",x"73",x"7c"),
   395 => (x"ff",x"c3",x"29",x"b7"),
   396 => (x"73",x"7c",x"71",x"99"),
   397 => (x"29",x"b7",x"d0",x"49"),
   398 => (x"71",x"99",x"ff",x"c3"),
   399 => (x"d8",x"49",x"73",x"7c"),
   400 => (x"7c",x"71",x"29",x"b7"),
   401 => (x"7c",x"7c",x"7c",x"c0"),
   402 => (x"7c",x"7c",x"7c",x"7c"),
   403 => (x"7c",x"7c",x"7c",x"7c"),
   404 => (x"78",x"e0",x"c0",x"7c"),
   405 => (x"dc",x"1e",x"66",x"c4"),
   406 => (x"d8",x"d2",x"ff",x"49"),
   407 => (x"73",x"86",x"c8",x"87"),
   408 => (x"ce",x"fa",x"26",x"48"),
   409 => (x"5b",x"5e",x"0e",x"87"),
   410 => (x"1e",x"0e",x"5d",x"5c"),
   411 => (x"d4",x"ff",x"7e",x"71"),
   412 => (x"c2",x"1e",x"6e",x"4b"),
   413 => (x"fe",x"49",x"de",x"f1"),
   414 => (x"c4",x"87",x"d2",x"c7"),
   415 => (x"9d",x"4d",x"70",x"86"),
   416 => (x"87",x"c3",x"c3",x"02"),
   417 => (x"bf",x"e6",x"f1",x"c2"),
   418 => (x"fe",x"49",x"6e",x"4c"),
   419 => (x"ff",x"87",x"f1",x"db"),
   420 => (x"c5",x"c8",x"48",x"d0"),
   421 => (x"7b",x"d6",x"c1",x"78"),
   422 => (x"7b",x"15",x"4a",x"c0"),
   423 => (x"e0",x"c0",x"82",x"c1"),
   424 => (x"f5",x"04",x"aa",x"b7"),
   425 => (x"48",x"d0",x"ff",x"87"),
   426 => (x"c5",x"c8",x"78",x"c4"),
   427 => (x"7b",x"d3",x"c1",x"78"),
   428 => (x"78",x"c4",x"7b",x"c1"),
   429 => (x"c1",x"02",x"9c",x"74"),
   430 => (x"df",x"c2",x"87",x"fc"),
   431 => (x"c0",x"c8",x"7e",x"e6"),
   432 => (x"b7",x"c0",x"8c",x"4d"),
   433 => (x"87",x"c6",x"03",x"ac"),
   434 => (x"4d",x"a4",x"c0",x"c8"),
   435 => (x"ec",x"c2",x"4c",x"c0"),
   436 => (x"49",x"bf",x"97",x"d7"),
   437 => (x"d2",x"02",x"99",x"d0"),
   438 => (x"c2",x"1e",x"c0",x"87"),
   439 => (x"fe",x"49",x"de",x"f1"),
   440 => (x"c4",x"87",x"c6",x"c9"),
   441 => (x"4a",x"49",x"70",x"86"),
   442 => (x"c2",x"87",x"ef",x"c0"),
   443 => (x"c2",x"1e",x"e6",x"df"),
   444 => (x"fe",x"49",x"de",x"f1"),
   445 => (x"c4",x"87",x"f2",x"c8"),
   446 => (x"4a",x"49",x"70",x"86"),
   447 => (x"c8",x"48",x"d0",x"ff"),
   448 => (x"d4",x"c1",x"78",x"c5"),
   449 => (x"bf",x"97",x"6e",x"7b"),
   450 => (x"c1",x"48",x"6e",x"7b"),
   451 => (x"c1",x"7e",x"70",x"80"),
   452 => (x"f0",x"ff",x"05",x"8d"),
   453 => (x"48",x"d0",x"ff",x"87"),
   454 => (x"9a",x"72",x"78",x"c4"),
   455 => (x"c0",x"87",x"c5",x"05"),
   456 => (x"87",x"e5",x"c0",x"48"),
   457 => (x"f1",x"c2",x"1e",x"c1"),
   458 => (x"c6",x"fe",x"49",x"de"),
   459 => (x"86",x"c4",x"87",x"da"),
   460 => (x"fe",x"05",x"9c",x"74"),
   461 => (x"d0",x"ff",x"87",x"c4"),
   462 => (x"78",x"c5",x"c8",x"48"),
   463 => (x"c0",x"7b",x"d3",x"c1"),
   464 => (x"c1",x"78",x"c4",x"7b"),
   465 => (x"c0",x"87",x"c2",x"48"),
   466 => (x"4d",x"26",x"26",x"48"),
   467 => (x"4b",x"26",x"4c",x"26"),
   468 => (x"5e",x"0e",x"4f",x"26"),
   469 => (x"71",x"0e",x"5c",x"5b"),
   470 => (x"02",x"66",x"cc",x"4b"),
   471 => (x"c0",x"4c",x"87",x"d8"),
   472 => (x"d8",x"02",x"8c",x"f0"),
   473 => (x"c1",x"4a",x"74",x"87"),
   474 => (x"87",x"d1",x"02",x"8a"),
   475 => (x"87",x"cd",x"02",x"8a"),
   476 => (x"87",x"c9",x"02",x"8a"),
   477 => (x"49",x"73",x"87",x"d7"),
   478 => (x"d0",x"87",x"ea",x"fb"),
   479 => (x"c0",x"1e",x"74",x"87"),
   480 => (x"87",x"e0",x"f9",x"49"),
   481 => (x"49",x"73",x"1e",x"74"),
   482 => (x"c8",x"87",x"d9",x"f9"),
   483 => (x"87",x"fc",x"fe",x"86"),
   484 => (x"de",x"c2",x"1e",x"00"),
   485 => (x"c1",x"49",x"bf",x"fa"),
   486 => (x"fe",x"de",x"c2",x"b9"),
   487 => (x"48",x"d4",x"ff",x"59"),
   488 => (x"ff",x"78",x"ff",x"c3"),
   489 => (x"e1",x"c8",x"48",x"d0"),
   490 => (x"48",x"d4",x"ff",x"78"),
   491 => (x"31",x"c4",x"78",x"c1"),
   492 => (x"d0",x"ff",x"78",x"71"),
   493 => (x"78",x"e0",x"c0",x"48"),
   494 => (x"00",x"00",x"4f",x"26"),
   495 => (x"00",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

