
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f4",x"f1",x"c2",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"f4",x"f1",x"c2"),
    14 => (x"48",x"c0",x"df",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"cd",x"dc"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"11",x"1e",x"4f"),
    50 => (x"78",x"08",x"d4",x"ff"),
    51 => (x"c1",x"48",x"66",x"c4"),
    52 => (x"58",x"a6",x"c8",x"88"),
    53 => (x"ed",x"05",x"98",x"70"),
    54 => (x"1e",x"4f",x"26",x"87"),
    55 => (x"c3",x"48",x"d4",x"ff"),
    56 => (x"51",x"68",x"78",x"ff"),
    57 => (x"c1",x"48",x"66",x"c4"),
    58 => (x"58",x"a6",x"c8",x"88"),
    59 => (x"eb",x"05",x"98",x"70"),
    60 => (x"1e",x"4f",x"26",x"87"),
    61 => (x"d4",x"ff",x"1e",x"73"),
    62 => (x"7b",x"ff",x"c3",x"4b"),
    63 => (x"ff",x"c3",x"4a",x"6b"),
    64 => (x"c8",x"49",x"6b",x"7b"),
    65 => (x"c3",x"b1",x"72",x"32"),
    66 => (x"4a",x"6b",x"7b",x"ff"),
    67 => (x"b2",x"71",x"31",x"c8"),
    68 => (x"6b",x"7b",x"ff",x"c3"),
    69 => (x"72",x"32",x"c8",x"49"),
    70 => (x"c4",x"48",x"71",x"b1"),
    71 => (x"26",x"4d",x"26",x"87"),
    72 => (x"26",x"4b",x"26",x"4c"),
    73 => (x"5b",x"5e",x"0e",x"4f"),
    74 => (x"71",x"0e",x"5d",x"5c"),
    75 => (x"4c",x"d4",x"ff",x"4a"),
    76 => (x"ff",x"c3",x"49",x"72"),
    77 => (x"c2",x"7c",x"71",x"99"),
    78 => (x"05",x"bf",x"c0",x"df"),
    79 => (x"66",x"d0",x"87",x"c8"),
    80 => (x"d4",x"30",x"c9",x"48"),
    81 => (x"66",x"d0",x"58",x"a6"),
    82 => (x"c3",x"29",x"d8",x"49"),
    83 => (x"7c",x"71",x"99",x"ff"),
    84 => (x"d0",x"49",x"66",x"d0"),
    85 => (x"99",x"ff",x"c3",x"29"),
    86 => (x"66",x"d0",x"7c",x"71"),
    87 => (x"c3",x"29",x"c8",x"49"),
    88 => (x"7c",x"71",x"99",x"ff"),
    89 => (x"c3",x"49",x"66",x"d0"),
    90 => (x"7c",x"71",x"99",x"ff"),
    91 => (x"29",x"d0",x"49",x"72"),
    92 => (x"71",x"99",x"ff",x"c3"),
    93 => (x"c9",x"4b",x"6c",x"7c"),
    94 => (x"c3",x"4d",x"ff",x"f0"),
    95 => (x"d0",x"05",x"ab",x"ff"),
    96 => (x"7c",x"ff",x"c3",x"87"),
    97 => (x"8d",x"c1",x"4b",x"6c"),
    98 => (x"c3",x"87",x"c6",x"02"),
    99 => (x"f0",x"02",x"ab",x"ff"),
   100 => (x"fe",x"48",x"73",x"87"),
   101 => (x"c0",x"1e",x"87",x"c7"),
   102 => (x"48",x"d4",x"ff",x"49"),
   103 => (x"c1",x"78",x"ff",x"c3"),
   104 => (x"b7",x"c8",x"c3",x"81"),
   105 => (x"87",x"f1",x"04",x"a9"),
   106 => (x"73",x"1e",x"4f",x"26"),
   107 => (x"c4",x"87",x"e7",x"1e"),
   108 => (x"c0",x"4b",x"df",x"f8"),
   109 => (x"f0",x"ff",x"c0",x"1e"),
   110 => (x"fd",x"49",x"f7",x"c1"),
   111 => (x"86",x"c4",x"87",x"e7"),
   112 => (x"c0",x"05",x"a8",x"c1"),
   113 => (x"d4",x"ff",x"87",x"ea"),
   114 => (x"78",x"ff",x"c3",x"48"),
   115 => (x"c0",x"c0",x"c0",x"c1"),
   116 => (x"c0",x"1e",x"c0",x"c0"),
   117 => (x"e9",x"c1",x"f0",x"e1"),
   118 => (x"87",x"c9",x"fd",x"49"),
   119 => (x"98",x"70",x"86",x"c4"),
   120 => (x"ff",x"87",x"ca",x"05"),
   121 => (x"ff",x"c3",x"48",x"d4"),
   122 => (x"cb",x"48",x"c1",x"78"),
   123 => (x"87",x"e6",x"fe",x"87"),
   124 => (x"fe",x"05",x"8b",x"c1"),
   125 => (x"48",x"c0",x"87",x"fd"),
   126 => (x"1e",x"87",x"e6",x"fc"),
   127 => (x"d4",x"ff",x"1e",x"73"),
   128 => (x"78",x"ff",x"c3",x"48"),
   129 => (x"1e",x"c0",x"4b",x"d3"),
   130 => (x"c1",x"f0",x"ff",x"c0"),
   131 => (x"d4",x"fc",x"49",x"c1"),
   132 => (x"70",x"86",x"c4",x"87"),
   133 => (x"87",x"ca",x"05",x"98"),
   134 => (x"c3",x"48",x"d4",x"ff"),
   135 => (x"48",x"c1",x"78",x"ff"),
   136 => (x"f1",x"fd",x"87",x"cb"),
   137 => (x"05",x"8b",x"c1",x"87"),
   138 => (x"c0",x"87",x"db",x"ff"),
   139 => (x"87",x"f1",x"fb",x"48"),
   140 => (x"5c",x"5b",x"5e",x"0e"),
   141 => (x"4c",x"d4",x"ff",x"0e"),
   142 => (x"c6",x"87",x"db",x"fd"),
   143 => (x"e1",x"c0",x"1e",x"ea"),
   144 => (x"49",x"c8",x"c1",x"f0"),
   145 => (x"c4",x"87",x"de",x"fb"),
   146 => (x"02",x"a8",x"c1",x"86"),
   147 => (x"ea",x"fe",x"87",x"c8"),
   148 => (x"c1",x"48",x"c0",x"87"),
   149 => (x"da",x"fa",x"87",x"e2"),
   150 => (x"cf",x"49",x"70",x"87"),
   151 => (x"c6",x"99",x"ff",x"ff"),
   152 => (x"c8",x"02",x"a9",x"ea"),
   153 => (x"87",x"d3",x"fe",x"87"),
   154 => (x"cb",x"c1",x"48",x"c0"),
   155 => (x"7c",x"ff",x"c3",x"87"),
   156 => (x"fc",x"4b",x"f1",x"c0"),
   157 => (x"98",x"70",x"87",x"f4"),
   158 => (x"87",x"eb",x"c0",x"02"),
   159 => (x"ff",x"c0",x"1e",x"c0"),
   160 => (x"49",x"fa",x"c1",x"f0"),
   161 => (x"c4",x"87",x"de",x"fa"),
   162 => (x"05",x"98",x"70",x"86"),
   163 => (x"ff",x"c3",x"87",x"d9"),
   164 => (x"c3",x"49",x"6c",x"7c"),
   165 => (x"7c",x"7c",x"7c",x"ff"),
   166 => (x"99",x"c0",x"c1",x"7c"),
   167 => (x"c1",x"87",x"c4",x"02"),
   168 => (x"c0",x"87",x"d5",x"48"),
   169 => (x"c2",x"87",x"d1",x"48"),
   170 => (x"87",x"c4",x"05",x"ab"),
   171 => (x"87",x"c8",x"48",x"c0"),
   172 => (x"fe",x"05",x"8b",x"c1"),
   173 => (x"48",x"c0",x"87",x"fd"),
   174 => (x"1e",x"87",x"e4",x"f9"),
   175 => (x"df",x"c2",x"1e",x"73"),
   176 => (x"78",x"c1",x"48",x"c0"),
   177 => (x"d0",x"ff",x"4b",x"c7"),
   178 => (x"fb",x"78",x"c2",x"48"),
   179 => (x"d0",x"ff",x"87",x"c8"),
   180 => (x"c0",x"78",x"c3",x"48"),
   181 => (x"d0",x"e5",x"c0",x"1e"),
   182 => (x"f9",x"49",x"c0",x"c1"),
   183 => (x"86",x"c4",x"87",x"c7"),
   184 => (x"c1",x"05",x"a8",x"c1"),
   185 => (x"ab",x"c2",x"4b",x"87"),
   186 => (x"c0",x"87",x"c5",x"05"),
   187 => (x"87",x"f9",x"c0",x"48"),
   188 => (x"ff",x"05",x"8b",x"c1"),
   189 => (x"f7",x"fc",x"87",x"d0"),
   190 => (x"c4",x"df",x"c2",x"87"),
   191 => (x"05",x"98",x"70",x"58"),
   192 => (x"1e",x"c1",x"87",x"cd"),
   193 => (x"c1",x"f0",x"ff",x"c0"),
   194 => (x"d8",x"f8",x"49",x"d0"),
   195 => (x"ff",x"86",x"c4",x"87"),
   196 => (x"ff",x"c3",x"48",x"d4"),
   197 => (x"87",x"e0",x"c4",x"78"),
   198 => (x"58",x"c8",x"df",x"c2"),
   199 => (x"c2",x"48",x"d0",x"ff"),
   200 => (x"48",x"d4",x"ff",x"78"),
   201 => (x"c1",x"78",x"ff",x"c3"),
   202 => (x"87",x"f5",x"f7",x"48"),
   203 => (x"5c",x"5b",x"5e",x"0e"),
   204 => (x"4a",x"71",x"0e",x"5d"),
   205 => (x"ff",x"4d",x"ff",x"c3"),
   206 => (x"7c",x"75",x"4c",x"d4"),
   207 => (x"c4",x"48",x"d0",x"ff"),
   208 => (x"7c",x"75",x"78",x"c3"),
   209 => (x"ff",x"c0",x"1e",x"72"),
   210 => (x"49",x"d8",x"c1",x"f0"),
   211 => (x"c4",x"87",x"d6",x"f7"),
   212 => (x"02",x"98",x"70",x"86"),
   213 => (x"48",x"c0",x"87",x"c5"),
   214 => (x"75",x"87",x"f0",x"c0"),
   215 => (x"7c",x"fe",x"c3",x"7c"),
   216 => (x"d4",x"1e",x"c0",x"c8"),
   217 => (x"dc",x"f5",x"49",x"66"),
   218 => (x"75",x"86",x"c4",x"87"),
   219 => (x"75",x"7c",x"75",x"7c"),
   220 => (x"e0",x"da",x"d8",x"7c"),
   221 => (x"6c",x"7c",x"75",x"4b"),
   222 => (x"c5",x"05",x"99",x"49"),
   223 => (x"05",x"8b",x"c1",x"87"),
   224 => (x"7c",x"75",x"87",x"f3"),
   225 => (x"c2",x"48",x"d0",x"ff"),
   226 => (x"f6",x"48",x"c1",x"78"),
   227 => (x"ff",x"1e",x"87",x"cf"),
   228 => (x"d0",x"ff",x"4a",x"d4"),
   229 => (x"78",x"d1",x"c4",x"48"),
   230 => (x"c1",x"7a",x"ff",x"c3"),
   231 => (x"87",x"f8",x"05",x"89"),
   232 => (x"73",x"1e",x"4f",x"26"),
   233 => (x"c5",x"4b",x"71",x"1e"),
   234 => (x"4a",x"df",x"cd",x"ee"),
   235 => (x"c3",x"48",x"d4",x"ff"),
   236 => (x"48",x"68",x"78",x"ff"),
   237 => (x"02",x"a8",x"fe",x"c3"),
   238 => (x"8a",x"c1",x"87",x"c5"),
   239 => (x"72",x"87",x"ed",x"05"),
   240 => (x"87",x"c5",x"05",x"9a"),
   241 => (x"ea",x"c0",x"48",x"c0"),
   242 => (x"02",x"9b",x"73",x"87"),
   243 => (x"66",x"c8",x"87",x"cc"),
   244 => (x"f4",x"49",x"73",x"1e"),
   245 => (x"86",x"c4",x"87",x"c5"),
   246 => (x"66",x"c8",x"87",x"c6"),
   247 => (x"87",x"ee",x"fe",x"49"),
   248 => (x"c3",x"48",x"d4",x"ff"),
   249 => (x"73",x"78",x"78",x"ff"),
   250 => (x"87",x"c5",x"05",x"9b"),
   251 => (x"d0",x"48",x"d0",x"ff"),
   252 => (x"f4",x"48",x"c1",x"78"),
   253 => (x"73",x"1e",x"87",x"eb"),
   254 => (x"c0",x"4a",x"71",x"1e"),
   255 => (x"48",x"d4",x"ff",x"4b"),
   256 => (x"ff",x"78",x"ff",x"c3"),
   257 => (x"c3",x"c4",x"48",x"d0"),
   258 => (x"48",x"d4",x"ff",x"78"),
   259 => (x"72",x"78",x"ff",x"c3"),
   260 => (x"f0",x"ff",x"c0",x"1e"),
   261 => (x"f4",x"49",x"d1",x"c1"),
   262 => (x"86",x"c4",x"87",x"cb"),
   263 => (x"cd",x"05",x"98",x"70"),
   264 => (x"1e",x"c0",x"c8",x"87"),
   265 => (x"fd",x"49",x"66",x"cc"),
   266 => (x"86",x"c4",x"87",x"f8"),
   267 => (x"d0",x"ff",x"4b",x"70"),
   268 => (x"73",x"78",x"c2",x"48"),
   269 => (x"87",x"e9",x"f3",x"48"),
   270 => (x"5c",x"5b",x"5e",x"0e"),
   271 => (x"1e",x"c0",x"0e",x"5d"),
   272 => (x"c1",x"f0",x"ff",x"c0"),
   273 => (x"dc",x"f3",x"49",x"c9"),
   274 => (x"c2",x"1e",x"d2",x"87"),
   275 => (x"fd",x"49",x"c8",x"df"),
   276 => (x"86",x"c8",x"87",x"d0"),
   277 => (x"84",x"c1",x"4c",x"c0"),
   278 => (x"04",x"ac",x"b7",x"d2"),
   279 => (x"df",x"c2",x"87",x"f8"),
   280 => (x"49",x"bf",x"97",x"c8"),
   281 => (x"c1",x"99",x"c0",x"c3"),
   282 => (x"c0",x"05",x"a9",x"c0"),
   283 => (x"df",x"c2",x"87",x"e7"),
   284 => (x"49",x"bf",x"97",x"cf"),
   285 => (x"df",x"c2",x"31",x"d0"),
   286 => (x"4a",x"bf",x"97",x"d0"),
   287 => (x"b1",x"72",x"32",x"c8"),
   288 => (x"97",x"d1",x"df",x"c2"),
   289 => (x"71",x"b1",x"4a",x"bf"),
   290 => (x"ff",x"ff",x"cf",x"4c"),
   291 => (x"84",x"c1",x"9c",x"ff"),
   292 => (x"e7",x"c1",x"34",x"ca"),
   293 => (x"d1",x"df",x"c2",x"87"),
   294 => (x"c1",x"49",x"bf",x"97"),
   295 => (x"c2",x"99",x"c6",x"31"),
   296 => (x"bf",x"97",x"d2",x"df"),
   297 => (x"2a",x"b7",x"c7",x"4a"),
   298 => (x"df",x"c2",x"b1",x"72"),
   299 => (x"4a",x"bf",x"97",x"cd"),
   300 => (x"c2",x"9d",x"cf",x"4d"),
   301 => (x"bf",x"97",x"ce",x"df"),
   302 => (x"ca",x"9a",x"c3",x"4a"),
   303 => (x"cf",x"df",x"c2",x"32"),
   304 => (x"c2",x"4b",x"bf",x"97"),
   305 => (x"c2",x"b2",x"73",x"33"),
   306 => (x"bf",x"97",x"d0",x"df"),
   307 => (x"9b",x"c0",x"c3",x"4b"),
   308 => (x"73",x"2b",x"b7",x"c6"),
   309 => (x"c1",x"81",x"c2",x"b2"),
   310 => (x"70",x"30",x"71",x"48"),
   311 => (x"75",x"48",x"c1",x"49"),
   312 => (x"72",x"4d",x"70",x"30"),
   313 => (x"71",x"84",x"c1",x"4c"),
   314 => (x"b7",x"c0",x"c8",x"94"),
   315 => (x"87",x"cc",x"06",x"ad"),
   316 => (x"2d",x"b7",x"34",x"c1"),
   317 => (x"ad",x"b7",x"c0",x"c8"),
   318 => (x"87",x"f4",x"ff",x"01"),
   319 => (x"dc",x"f0",x"48",x"74"),
   320 => (x"5b",x"5e",x"0e",x"87"),
   321 => (x"f8",x"0e",x"5d",x"5c"),
   322 => (x"ee",x"e7",x"c2",x"86"),
   323 => (x"c2",x"78",x"c0",x"48"),
   324 => (x"c0",x"1e",x"e6",x"df"),
   325 => (x"87",x"de",x"fb",x"49"),
   326 => (x"98",x"70",x"86",x"c4"),
   327 => (x"c0",x"87",x"c5",x"05"),
   328 => (x"87",x"ce",x"c9",x"48"),
   329 => (x"7e",x"c1",x"4d",x"c0"),
   330 => (x"bf",x"cb",x"f2",x"c0"),
   331 => (x"dc",x"e0",x"c2",x"49"),
   332 => (x"4b",x"c8",x"71",x"4a"),
   333 => (x"70",x"87",x"f3",x"ec"),
   334 => (x"87",x"c2",x"05",x"98"),
   335 => (x"f2",x"c0",x"7e",x"c0"),
   336 => (x"c2",x"49",x"bf",x"c7"),
   337 => (x"71",x"4a",x"f8",x"e0"),
   338 => (x"dd",x"ec",x"4b",x"c8"),
   339 => (x"05",x"98",x"70",x"87"),
   340 => (x"7e",x"c0",x"87",x"c2"),
   341 => (x"fd",x"c0",x"02",x"6e"),
   342 => (x"ec",x"e6",x"c2",x"87"),
   343 => (x"e7",x"c2",x"4d",x"bf"),
   344 => (x"7e",x"bf",x"9f",x"e4"),
   345 => (x"ea",x"d6",x"c5",x"48"),
   346 => (x"87",x"c7",x"05",x"a8"),
   347 => (x"bf",x"ec",x"e6",x"c2"),
   348 => (x"6e",x"87",x"ce",x"4d"),
   349 => (x"d5",x"e9",x"ca",x"48"),
   350 => (x"87",x"c5",x"02",x"a8"),
   351 => (x"f1",x"c7",x"48",x"c0"),
   352 => (x"e6",x"df",x"c2",x"87"),
   353 => (x"f9",x"49",x"75",x"1e"),
   354 => (x"86",x"c4",x"87",x"ec"),
   355 => (x"c5",x"05",x"98",x"70"),
   356 => (x"c7",x"48",x"c0",x"87"),
   357 => (x"f2",x"c0",x"87",x"dc"),
   358 => (x"c2",x"49",x"bf",x"c7"),
   359 => (x"71",x"4a",x"f8",x"e0"),
   360 => (x"c5",x"eb",x"4b",x"c8"),
   361 => (x"05",x"98",x"70",x"87"),
   362 => (x"e7",x"c2",x"87",x"c8"),
   363 => (x"78",x"c1",x"48",x"ee"),
   364 => (x"f2",x"c0",x"87",x"da"),
   365 => (x"c2",x"49",x"bf",x"cb"),
   366 => (x"71",x"4a",x"dc",x"e0"),
   367 => (x"e9",x"ea",x"4b",x"c8"),
   368 => (x"02",x"98",x"70",x"87"),
   369 => (x"c0",x"87",x"c5",x"c0"),
   370 => (x"87",x"e6",x"c6",x"48"),
   371 => (x"97",x"e4",x"e7",x"c2"),
   372 => (x"d5",x"c1",x"49",x"bf"),
   373 => (x"cd",x"c0",x"05",x"a9"),
   374 => (x"e5",x"e7",x"c2",x"87"),
   375 => (x"c2",x"49",x"bf",x"97"),
   376 => (x"c0",x"02",x"a9",x"ea"),
   377 => (x"48",x"c0",x"87",x"c5"),
   378 => (x"c2",x"87",x"c7",x"c6"),
   379 => (x"bf",x"97",x"e6",x"df"),
   380 => (x"e9",x"c3",x"48",x"7e"),
   381 => (x"ce",x"c0",x"02",x"a8"),
   382 => (x"c3",x"48",x"6e",x"87"),
   383 => (x"c0",x"02",x"a8",x"eb"),
   384 => (x"48",x"c0",x"87",x"c5"),
   385 => (x"c2",x"87",x"eb",x"c5"),
   386 => (x"bf",x"97",x"f1",x"df"),
   387 => (x"c0",x"05",x"99",x"49"),
   388 => (x"df",x"c2",x"87",x"cc"),
   389 => (x"49",x"bf",x"97",x"f2"),
   390 => (x"c0",x"02",x"a9",x"c2"),
   391 => (x"48",x"c0",x"87",x"c5"),
   392 => (x"c2",x"87",x"cf",x"c5"),
   393 => (x"bf",x"97",x"f3",x"df"),
   394 => (x"ea",x"e7",x"c2",x"48"),
   395 => (x"48",x"4c",x"70",x"58"),
   396 => (x"e7",x"c2",x"88",x"c1"),
   397 => (x"df",x"c2",x"58",x"ee"),
   398 => (x"49",x"bf",x"97",x"f4"),
   399 => (x"df",x"c2",x"81",x"75"),
   400 => (x"4a",x"bf",x"97",x"f5"),
   401 => (x"a1",x"72",x"32",x"c8"),
   402 => (x"fb",x"eb",x"c2",x"7e"),
   403 => (x"c2",x"78",x"6e",x"48"),
   404 => (x"bf",x"97",x"f6",x"df"),
   405 => (x"58",x"a6",x"c8",x"48"),
   406 => (x"bf",x"ee",x"e7",x"c2"),
   407 => (x"87",x"d4",x"c2",x"02"),
   408 => (x"bf",x"c7",x"f2",x"c0"),
   409 => (x"f8",x"e0",x"c2",x"49"),
   410 => (x"4b",x"c8",x"71",x"4a"),
   411 => (x"70",x"87",x"fb",x"e7"),
   412 => (x"c5",x"c0",x"02",x"98"),
   413 => (x"c3",x"48",x"c0",x"87"),
   414 => (x"e7",x"c2",x"87",x"f8"),
   415 => (x"c2",x"4c",x"bf",x"e6"),
   416 => (x"c2",x"5c",x"cf",x"ec"),
   417 => (x"bf",x"97",x"cb",x"e0"),
   418 => (x"c2",x"31",x"c8",x"49"),
   419 => (x"bf",x"97",x"ca",x"e0"),
   420 => (x"c2",x"49",x"a1",x"4a"),
   421 => (x"bf",x"97",x"cc",x"e0"),
   422 => (x"72",x"32",x"d0",x"4a"),
   423 => (x"e0",x"c2",x"49",x"a1"),
   424 => (x"4a",x"bf",x"97",x"cd"),
   425 => (x"a1",x"72",x"32",x"d8"),
   426 => (x"91",x"66",x"c4",x"49"),
   427 => (x"bf",x"fb",x"eb",x"c2"),
   428 => (x"c3",x"ec",x"c2",x"81"),
   429 => (x"d3",x"e0",x"c2",x"59"),
   430 => (x"c8",x"4a",x"bf",x"97"),
   431 => (x"d2",x"e0",x"c2",x"32"),
   432 => (x"a2",x"4b",x"bf",x"97"),
   433 => (x"d4",x"e0",x"c2",x"4a"),
   434 => (x"d0",x"4b",x"bf",x"97"),
   435 => (x"4a",x"a2",x"73",x"33"),
   436 => (x"97",x"d5",x"e0",x"c2"),
   437 => (x"9b",x"cf",x"4b",x"bf"),
   438 => (x"a2",x"73",x"33",x"d8"),
   439 => (x"c7",x"ec",x"c2",x"4a"),
   440 => (x"c3",x"ec",x"c2",x"5a"),
   441 => (x"8a",x"c2",x"4a",x"bf"),
   442 => (x"ec",x"c2",x"92",x"74"),
   443 => (x"a1",x"72",x"48",x"c7"),
   444 => (x"87",x"ca",x"c1",x"78"),
   445 => (x"97",x"f8",x"df",x"c2"),
   446 => (x"31",x"c8",x"49",x"bf"),
   447 => (x"97",x"f7",x"df",x"c2"),
   448 => (x"49",x"a1",x"4a",x"bf"),
   449 => (x"59",x"f6",x"e7",x"c2"),
   450 => (x"bf",x"f2",x"e7",x"c2"),
   451 => (x"c7",x"31",x"c5",x"49"),
   452 => (x"29",x"c9",x"81",x"ff"),
   453 => (x"59",x"cf",x"ec",x"c2"),
   454 => (x"97",x"fd",x"df",x"c2"),
   455 => (x"32",x"c8",x"4a",x"bf"),
   456 => (x"97",x"fc",x"df",x"c2"),
   457 => (x"4a",x"a2",x"4b",x"bf"),
   458 => (x"6e",x"92",x"66",x"c4"),
   459 => (x"cb",x"ec",x"c2",x"82"),
   460 => (x"c3",x"ec",x"c2",x"5a"),
   461 => (x"c2",x"78",x"c0",x"48"),
   462 => (x"72",x"48",x"ff",x"eb"),
   463 => (x"ec",x"c2",x"78",x"a1"),
   464 => (x"ec",x"c2",x"48",x"cf"),
   465 => (x"c2",x"78",x"bf",x"c3"),
   466 => (x"c2",x"48",x"d3",x"ec"),
   467 => (x"78",x"bf",x"c7",x"ec"),
   468 => (x"bf",x"ee",x"e7",x"c2"),
   469 => (x"87",x"c9",x"c0",x"02"),
   470 => (x"30",x"c4",x"48",x"74"),
   471 => (x"c9",x"c0",x"7e",x"70"),
   472 => (x"cb",x"ec",x"c2",x"87"),
   473 => (x"30",x"c4",x"48",x"bf"),
   474 => (x"e7",x"c2",x"7e",x"70"),
   475 => (x"78",x"6e",x"48",x"f2"),
   476 => (x"8e",x"f8",x"48",x"c1"),
   477 => (x"4c",x"26",x"4d",x"26"),
   478 => (x"4f",x"26",x"4b",x"26"),
   479 => (x"5c",x"5b",x"5e",x"0e"),
   480 => (x"4a",x"71",x"0e",x"5d"),
   481 => (x"bf",x"ee",x"e7",x"c2"),
   482 => (x"72",x"87",x"cb",x"02"),
   483 => (x"72",x"2b",x"c7",x"4b"),
   484 => (x"9c",x"ff",x"c1",x"4c"),
   485 => (x"4b",x"72",x"87",x"c9"),
   486 => (x"4c",x"72",x"2b",x"c8"),
   487 => (x"c2",x"9c",x"ff",x"c3"),
   488 => (x"83",x"bf",x"fb",x"eb"),
   489 => (x"bf",x"c3",x"f2",x"c0"),
   490 => (x"87",x"d9",x"02",x"ab"),
   491 => (x"5b",x"c7",x"f2",x"c0"),
   492 => (x"1e",x"e6",x"df",x"c2"),
   493 => (x"fd",x"f0",x"49",x"73"),
   494 => (x"70",x"86",x"c4",x"87"),
   495 => (x"87",x"c5",x"05",x"98"),
   496 => (x"e6",x"c0",x"48",x"c0"),
   497 => (x"ee",x"e7",x"c2",x"87"),
   498 => (x"87",x"d2",x"02",x"bf"),
   499 => (x"91",x"c4",x"49",x"74"),
   500 => (x"81",x"e6",x"df",x"c2"),
   501 => (x"ff",x"cf",x"4d",x"69"),
   502 => (x"9d",x"ff",x"ff",x"ff"),
   503 => (x"49",x"74",x"87",x"cb"),
   504 => (x"df",x"c2",x"91",x"c2"),
   505 => (x"69",x"9f",x"81",x"e6"),
   506 => (x"fe",x"48",x"75",x"4d"),
   507 => (x"5e",x"0e",x"87",x"c6"),
   508 => (x"0e",x"5d",x"5c",x"5b"),
   509 => (x"c0",x"4d",x"71",x"1e"),
   510 => (x"ca",x"49",x"c1",x"1e"),
   511 => (x"86",x"c4",x"87",x"ee"),
   512 => (x"02",x"9c",x"4c",x"70"),
   513 => (x"c2",x"87",x"c0",x"c1"),
   514 => (x"75",x"4a",x"f6",x"e7"),
   515 => (x"87",x"ff",x"e0",x"49"),
   516 => (x"c0",x"02",x"98",x"70"),
   517 => (x"4a",x"74",x"87",x"f1"),
   518 => (x"4b",x"cb",x"49",x"75"),
   519 => (x"70",x"87",x"e5",x"e1"),
   520 => (x"e2",x"c0",x"02",x"98"),
   521 => (x"74",x"1e",x"c0",x"87"),
   522 => (x"87",x"c7",x"02",x"9c"),
   523 => (x"c0",x"48",x"a6",x"c4"),
   524 => (x"c4",x"87",x"c5",x"78"),
   525 => (x"78",x"c1",x"48",x"a6"),
   526 => (x"c9",x"49",x"66",x"c4"),
   527 => (x"86",x"c4",x"87",x"ee"),
   528 => (x"05",x"9c",x"4c",x"70"),
   529 => (x"74",x"87",x"c0",x"ff"),
   530 => (x"e7",x"fc",x"26",x"48"),
   531 => (x"5b",x"5e",x"0e",x"87"),
   532 => (x"1e",x"0e",x"5d",x"5c"),
   533 => (x"05",x"9b",x"4b",x"71"),
   534 => (x"48",x"c0",x"87",x"c5"),
   535 => (x"c8",x"87",x"e5",x"c1"),
   536 => (x"7d",x"c0",x"4d",x"a3"),
   537 => (x"c7",x"02",x"66",x"d4"),
   538 => (x"97",x"66",x"d4",x"87"),
   539 => (x"87",x"c5",x"05",x"bf"),
   540 => (x"cf",x"c1",x"48",x"c0"),
   541 => (x"49",x"66",x"d4",x"87"),
   542 => (x"70",x"87",x"f3",x"fd"),
   543 => (x"c1",x"02",x"9c",x"4c"),
   544 => (x"a4",x"dc",x"87",x"c0"),
   545 => (x"da",x"7d",x"69",x"49"),
   546 => (x"a3",x"c4",x"49",x"a4"),
   547 => (x"7a",x"69",x"9f",x"4a"),
   548 => (x"bf",x"ee",x"e7",x"c2"),
   549 => (x"d4",x"87",x"d2",x"02"),
   550 => (x"69",x"9f",x"49",x"a4"),
   551 => (x"ff",x"ff",x"c0",x"49"),
   552 => (x"d0",x"48",x"71",x"99"),
   553 => (x"c2",x"7e",x"70",x"30"),
   554 => (x"6e",x"7e",x"c0",x"87"),
   555 => (x"80",x"6a",x"48",x"49"),
   556 => (x"7b",x"c0",x"7a",x"70"),
   557 => (x"6a",x"49",x"a3",x"cc"),
   558 => (x"49",x"a3",x"d0",x"79"),
   559 => (x"48",x"74",x"79",x"c0"),
   560 => (x"48",x"c0",x"87",x"c2"),
   561 => (x"87",x"ec",x"fa",x"26"),
   562 => (x"5c",x"5b",x"5e",x"0e"),
   563 => (x"4c",x"71",x"0e",x"5d"),
   564 => (x"48",x"c3",x"f2",x"c0"),
   565 => (x"9c",x"74",x"78",x"ff"),
   566 => (x"87",x"ca",x"c1",x"02"),
   567 => (x"69",x"49",x"a4",x"c8"),
   568 => (x"87",x"c2",x"c1",x"02"),
   569 => (x"6c",x"4a",x"66",x"d0"),
   570 => (x"a6",x"d4",x"82",x"49"),
   571 => (x"4d",x"66",x"d0",x"5a"),
   572 => (x"ea",x"e7",x"c2",x"b9"),
   573 => (x"ba",x"ff",x"4a",x"bf"),
   574 => (x"99",x"71",x"99",x"72"),
   575 => (x"87",x"e4",x"c0",x"02"),
   576 => (x"6b",x"4b",x"a4",x"c4"),
   577 => (x"87",x"f4",x"f9",x"49"),
   578 => (x"e7",x"c2",x"7b",x"70"),
   579 => (x"6c",x"49",x"bf",x"e6"),
   580 => (x"75",x"7c",x"71",x"81"),
   581 => (x"ea",x"e7",x"c2",x"b9"),
   582 => (x"ba",x"ff",x"4a",x"bf"),
   583 => (x"99",x"71",x"99",x"72"),
   584 => (x"87",x"dc",x"ff",x"05"),
   585 => (x"cb",x"f9",x"7c",x"75"),
   586 => (x"1e",x"73",x"1e",x"87"),
   587 => (x"02",x"9b",x"4b",x"71"),
   588 => (x"a3",x"c8",x"87",x"c7"),
   589 => (x"c5",x"05",x"69",x"49"),
   590 => (x"c0",x"48",x"c0",x"87"),
   591 => (x"eb",x"c2",x"87",x"eb"),
   592 => (x"c4",x"4a",x"bf",x"ff"),
   593 => (x"49",x"69",x"49",x"a3"),
   594 => (x"e7",x"c2",x"89",x"c2"),
   595 => (x"71",x"91",x"bf",x"e6"),
   596 => (x"e7",x"c2",x"4a",x"a2"),
   597 => (x"6b",x"49",x"bf",x"ea"),
   598 => (x"4a",x"a2",x"71",x"99"),
   599 => (x"72",x"1e",x"66",x"c8"),
   600 => (x"87",x"d2",x"ea",x"49"),
   601 => (x"49",x"70",x"86",x"c4"),
   602 => (x"87",x"cc",x"f8",x"48"),
   603 => (x"71",x"1e",x"73",x"1e"),
   604 => (x"c7",x"02",x"9b",x"4b"),
   605 => (x"49",x"a3",x"c8",x"87"),
   606 => (x"87",x"c5",x"05",x"69"),
   607 => (x"eb",x"c0",x"48",x"c0"),
   608 => (x"ff",x"eb",x"c2",x"87"),
   609 => (x"a3",x"c4",x"4a",x"bf"),
   610 => (x"c2",x"49",x"69",x"49"),
   611 => (x"e6",x"e7",x"c2",x"89"),
   612 => (x"a2",x"71",x"91",x"bf"),
   613 => (x"ea",x"e7",x"c2",x"4a"),
   614 => (x"99",x"6b",x"49",x"bf"),
   615 => (x"c8",x"4a",x"a2",x"71"),
   616 => (x"49",x"72",x"1e",x"66"),
   617 => (x"c4",x"87",x"c5",x"e6"),
   618 => (x"48",x"49",x"70",x"86"),
   619 => (x"0e",x"87",x"c9",x"f7"),
   620 => (x"5d",x"5c",x"5b",x"5e"),
   621 => (x"4b",x"71",x"1e",x"0e"),
   622 => (x"c9",x"4c",x"66",x"d4"),
   623 => (x"02",x"9b",x"73",x"2c"),
   624 => (x"c8",x"87",x"cf",x"c1"),
   625 => (x"02",x"69",x"49",x"a3"),
   626 => (x"d0",x"87",x"c7",x"c1"),
   627 => (x"66",x"d4",x"4d",x"a3"),
   628 => (x"ea",x"e7",x"c2",x"7d"),
   629 => (x"b9",x"ff",x"49",x"bf"),
   630 => (x"7e",x"99",x"4a",x"6b"),
   631 => (x"cd",x"03",x"ac",x"71"),
   632 => (x"7d",x"7b",x"c0",x"87"),
   633 => (x"c4",x"4a",x"a3",x"cc"),
   634 => (x"79",x"6a",x"49",x"a3"),
   635 => (x"8c",x"72",x"87",x"c2"),
   636 => (x"dd",x"02",x"9c",x"74"),
   637 => (x"73",x"1e",x"49",x"87"),
   638 => (x"87",x"cc",x"fb",x"49"),
   639 => (x"66",x"d4",x"86",x"c4"),
   640 => (x"99",x"ff",x"c7",x"49"),
   641 => (x"c2",x"87",x"cb",x"02"),
   642 => (x"73",x"1e",x"e6",x"df"),
   643 => (x"87",x"d9",x"fc",x"49"),
   644 => (x"f5",x"26",x"86",x"c4"),
   645 => (x"73",x"1e",x"87",x"de"),
   646 => (x"9b",x"4b",x"71",x"1e"),
   647 => (x"87",x"e4",x"c0",x"02"),
   648 => (x"5b",x"d3",x"ec",x"c2"),
   649 => (x"8a",x"c2",x"4a",x"73"),
   650 => (x"bf",x"e6",x"e7",x"c2"),
   651 => (x"eb",x"c2",x"92",x"49"),
   652 => (x"72",x"48",x"bf",x"ff"),
   653 => (x"d7",x"ec",x"c2",x"80"),
   654 => (x"c4",x"48",x"71",x"58"),
   655 => (x"f6",x"e7",x"c2",x"30"),
   656 => (x"87",x"ed",x"c0",x"58"),
   657 => (x"48",x"cf",x"ec",x"c2"),
   658 => (x"bf",x"c3",x"ec",x"c2"),
   659 => (x"d3",x"ec",x"c2",x"78"),
   660 => (x"c7",x"ec",x"c2",x"48"),
   661 => (x"e7",x"c2",x"78",x"bf"),
   662 => (x"c9",x"02",x"bf",x"ee"),
   663 => (x"e6",x"e7",x"c2",x"87"),
   664 => (x"31",x"c4",x"49",x"bf"),
   665 => (x"ec",x"c2",x"87",x"c7"),
   666 => (x"c4",x"49",x"bf",x"cb"),
   667 => (x"f6",x"e7",x"c2",x"31"),
   668 => (x"87",x"c4",x"f4",x"59"),
   669 => (x"5c",x"5b",x"5e",x"0e"),
   670 => (x"c0",x"4a",x"71",x"0e"),
   671 => (x"02",x"9a",x"72",x"4b"),
   672 => (x"da",x"87",x"e1",x"c0"),
   673 => (x"69",x"9f",x"49",x"a2"),
   674 => (x"ee",x"e7",x"c2",x"4b"),
   675 => (x"87",x"cf",x"02",x"bf"),
   676 => (x"9f",x"49",x"a2",x"d4"),
   677 => (x"c0",x"4c",x"49",x"69"),
   678 => (x"d0",x"9c",x"ff",x"ff"),
   679 => (x"c0",x"87",x"c2",x"34"),
   680 => (x"b3",x"49",x"74",x"4c"),
   681 => (x"ed",x"fd",x"49",x"73"),
   682 => (x"87",x"ca",x"f3",x"87"),
   683 => (x"5c",x"5b",x"5e",x"0e"),
   684 => (x"86",x"f4",x"0e",x"5d"),
   685 => (x"7e",x"c0",x"4a",x"71"),
   686 => (x"d8",x"02",x"9a",x"72"),
   687 => (x"e2",x"df",x"c2",x"87"),
   688 => (x"c2",x"78",x"c0",x"48"),
   689 => (x"c2",x"48",x"da",x"df"),
   690 => (x"78",x"bf",x"d3",x"ec"),
   691 => (x"48",x"de",x"df",x"c2"),
   692 => (x"bf",x"cf",x"ec",x"c2"),
   693 => (x"c3",x"e8",x"c2",x"78"),
   694 => (x"c2",x"50",x"c0",x"48"),
   695 => (x"49",x"bf",x"f2",x"e7"),
   696 => (x"bf",x"e2",x"df",x"c2"),
   697 => (x"03",x"aa",x"71",x"4a"),
   698 => (x"72",x"87",x"ff",x"c3"),
   699 => (x"05",x"99",x"cf",x"49"),
   700 => (x"c2",x"87",x"e0",x"c0"),
   701 => (x"c2",x"1e",x"e6",x"df"),
   702 => (x"49",x"bf",x"da",x"df"),
   703 => (x"48",x"da",x"df",x"c2"),
   704 => (x"71",x"78",x"a1",x"c1"),
   705 => (x"c4",x"87",x"ef",x"e3"),
   706 => (x"ff",x"f1",x"c0",x"86"),
   707 => (x"e6",x"df",x"c2",x"48"),
   708 => (x"c0",x"87",x"cc",x"78"),
   709 => (x"48",x"bf",x"ff",x"f1"),
   710 => (x"c0",x"80",x"e0",x"c0"),
   711 => (x"c2",x"58",x"c3",x"f2"),
   712 => (x"48",x"bf",x"e2",x"df"),
   713 => (x"df",x"c2",x"80",x"c1"),
   714 => (x"7f",x"27",x"58",x"e6"),
   715 => (x"bf",x"00",x"00",x"0c"),
   716 => (x"9d",x"4d",x"bf",x"97"),
   717 => (x"87",x"e2",x"c2",x"02"),
   718 => (x"02",x"ad",x"e5",x"c3"),
   719 => (x"c0",x"87",x"db",x"c2"),
   720 => (x"4b",x"bf",x"ff",x"f1"),
   721 => (x"11",x"49",x"a3",x"cb"),
   722 => (x"05",x"ac",x"cf",x"4c"),
   723 => (x"75",x"87",x"d2",x"c1"),
   724 => (x"c1",x"99",x"df",x"49"),
   725 => (x"c2",x"91",x"cd",x"89"),
   726 => (x"c1",x"81",x"f6",x"e7"),
   727 => (x"51",x"12",x"4a",x"a3"),
   728 => (x"12",x"4a",x"a3",x"c3"),
   729 => (x"4a",x"a3",x"c5",x"51"),
   730 => (x"a3",x"c7",x"51",x"12"),
   731 => (x"c9",x"51",x"12",x"4a"),
   732 => (x"51",x"12",x"4a",x"a3"),
   733 => (x"12",x"4a",x"a3",x"ce"),
   734 => (x"4a",x"a3",x"d0",x"51"),
   735 => (x"a3",x"d2",x"51",x"12"),
   736 => (x"d4",x"51",x"12",x"4a"),
   737 => (x"51",x"12",x"4a",x"a3"),
   738 => (x"12",x"4a",x"a3",x"d6"),
   739 => (x"4a",x"a3",x"d8",x"51"),
   740 => (x"a3",x"dc",x"51",x"12"),
   741 => (x"de",x"51",x"12",x"4a"),
   742 => (x"51",x"12",x"4a",x"a3"),
   743 => (x"f9",x"c0",x"7e",x"c1"),
   744 => (x"c8",x"49",x"74",x"87"),
   745 => (x"ea",x"c0",x"05",x"99"),
   746 => (x"d0",x"49",x"74",x"87"),
   747 => (x"87",x"d0",x"05",x"99"),
   748 => (x"c0",x"02",x"66",x"dc"),
   749 => (x"49",x"73",x"87",x"ca"),
   750 => (x"70",x"0f",x"66",x"dc"),
   751 => (x"87",x"d3",x"02",x"98"),
   752 => (x"c6",x"c0",x"05",x"6e"),
   753 => (x"f6",x"e7",x"c2",x"87"),
   754 => (x"c0",x"50",x"c0",x"48"),
   755 => (x"48",x"bf",x"ff",x"f1"),
   756 => (x"c2",x"87",x"e7",x"c2"),
   757 => (x"c0",x"48",x"c3",x"e8"),
   758 => (x"e7",x"c2",x"7e",x"50"),
   759 => (x"c2",x"49",x"bf",x"f2"),
   760 => (x"4a",x"bf",x"e2",x"df"),
   761 => (x"fc",x"04",x"aa",x"71"),
   762 => (x"ec",x"c2",x"87",x"c1"),
   763 => (x"c0",x"05",x"bf",x"d3"),
   764 => (x"e7",x"c2",x"87",x"c8"),
   765 => (x"c1",x"02",x"bf",x"ee"),
   766 => (x"f2",x"c0",x"87",x"fe"),
   767 => (x"78",x"ff",x"48",x"c3"),
   768 => (x"bf",x"de",x"df",x"c2"),
   769 => (x"87",x"f4",x"ed",x"49"),
   770 => (x"df",x"c2",x"49",x"70"),
   771 => (x"a6",x"c4",x"59",x"e2"),
   772 => (x"de",x"df",x"c2",x"48"),
   773 => (x"e7",x"c2",x"78",x"bf"),
   774 => (x"c0",x"02",x"bf",x"ee"),
   775 => (x"66",x"c4",x"87",x"d8"),
   776 => (x"ff",x"ff",x"cf",x"49"),
   777 => (x"a9",x"99",x"f8",x"ff"),
   778 => (x"87",x"c5",x"c0",x"02"),
   779 => (x"e1",x"c0",x"4d",x"c0"),
   780 => (x"c0",x"4d",x"c1",x"87"),
   781 => (x"66",x"c4",x"87",x"dc"),
   782 => (x"f8",x"ff",x"cf",x"49"),
   783 => (x"c0",x"02",x"a9",x"99"),
   784 => (x"a6",x"c8",x"87",x"c8"),
   785 => (x"c0",x"78",x"c0",x"48"),
   786 => (x"a6",x"c8",x"87",x"c5"),
   787 => (x"c8",x"78",x"c1",x"48"),
   788 => (x"9d",x"75",x"4d",x"66"),
   789 => (x"87",x"e0",x"c0",x"05"),
   790 => (x"c2",x"49",x"66",x"c4"),
   791 => (x"e6",x"e7",x"c2",x"89"),
   792 => (x"c2",x"91",x"4a",x"bf"),
   793 => (x"4a",x"bf",x"ff",x"eb"),
   794 => (x"48",x"da",x"df",x"c2"),
   795 => (x"c2",x"78",x"a1",x"72"),
   796 => (x"c0",x"48",x"e2",x"df"),
   797 => (x"87",x"e3",x"f9",x"78"),
   798 => (x"8e",x"f4",x"48",x"c0"),
   799 => (x"00",x"87",x"f5",x"eb"),
   800 => (x"ff",x"00",x"00",x"00"),
   801 => (x"8f",x"ff",x"ff",x"ff"),
   802 => (x"98",x"00",x"00",x"0c"),
   803 => (x"46",x"00",x"00",x"0c"),
   804 => (x"32",x"33",x"54",x"41"),
   805 => (x"00",x"20",x"20",x"20"),
   806 => (x"31",x"54",x"41",x"46"),
   807 => (x"20",x"20",x"20",x"36"),
   808 => (x"d4",x"ff",x"1e",x"00"),
   809 => (x"78",x"ff",x"c3",x"48"),
   810 => (x"4f",x"26",x"48",x"68"),
   811 => (x"48",x"d4",x"ff",x"1e"),
   812 => (x"ff",x"78",x"ff",x"c3"),
   813 => (x"e1",x"c8",x"48",x"d0"),
   814 => (x"48",x"d4",x"ff",x"78"),
   815 => (x"ec",x"c2",x"78",x"d4"),
   816 => (x"d4",x"ff",x"48",x"d7"),
   817 => (x"4f",x"26",x"50",x"bf"),
   818 => (x"48",x"d0",x"ff",x"1e"),
   819 => (x"26",x"78",x"e0",x"c0"),
   820 => (x"cc",x"ff",x"1e",x"4f"),
   821 => (x"99",x"49",x"70",x"87"),
   822 => (x"c0",x"87",x"c6",x"02"),
   823 => (x"f1",x"05",x"a9",x"fb"),
   824 => (x"26",x"48",x"71",x"87"),
   825 => (x"5b",x"5e",x"0e",x"4f"),
   826 => (x"4b",x"71",x"0e",x"5c"),
   827 => (x"f0",x"fe",x"4c",x"c0"),
   828 => (x"99",x"49",x"70",x"87"),
   829 => (x"87",x"f9",x"c0",x"02"),
   830 => (x"02",x"a9",x"ec",x"c0"),
   831 => (x"c0",x"87",x"f2",x"c0"),
   832 => (x"c0",x"02",x"a9",x"fb"),
   833 => (x"66",x"cc",x"87",x"eb"),
   834 => (x"c7",x"03",x"ac",x"b7"),
   835 => (x"02",x"66",x"d0",x"87"),
   836 => (x"53",x"71",x"87",x"c2"),
   837 => (x"c2",x"02",x"99",x"71"),
   838 => (x"fe",x"84",x"c1",x"87"),
   839 => (x"49",x"70",x"87",x"c3"),
   840 => (x"87",x"cd",x"02",x"99"),
   841 => (x"02",x"a9",x"ec",x"c0"),
   842 => (x"fb",x"c0",x"87",x"c7"),
   843 => (x"d5",x"ff",x"05",x"a9"),
   844 => (x"02",x"66",x"d0",x"87"),
   845 => (x"97",x"c0",x"87",x"c3"),
   846 => (x"a9",x"ec",x"c0",x"7b"),
   847 => (x"74",x"87",x"c4",x"05"),
   848 => (x"74",x"87",x"c5",x"4a"),
   849 => (x"8a",x"0a",x"c0",x"4a"),
   850 => (x"87",x"c2",x"48",x"72"),
   851 => (x"4c",x"26",x"4d",x"26"),
   852 => (x"4f",x"26",x"4b",x"26"),
   853 => (x"87",x"c9",x"fd",x"1e"),
   854 => (x"f0",x"c0",x"49",x"70"),
   855 => (x"ca",x"04",x"a9",x"b7"),
   856 => (x"b7",x"f9",x"c0",x"87"),
   857 => (x"87",x"c3",x"01",x"a9"),
   858 => (x"c1",x"89",x"f0",x"c0"),
   859 => (x"04",x"a9",x"b7",x"c1"),
   860 => (x"da",x"c1",x"87",x"ca"),
   861 => (x"c3",x"01",x"a9",x"b7"),
   862 => (x"89",x"f7",x"c0",x"87"),
   863 => (x"4f",x"26",x"48",x"71"),
   864 => (x"5c",x"5b",x"5e",x"0e"),
   865 => (x"ff",x"4a",x"71",x"0e"),
   866 => (x"49",x"72",x"4c",x"d4"),
   867 => (x"70",x"87",x"ea",x"c0"),
   868 => (x"c2",x"02",x"9b",x"4b"),
   869 => (x"ff",x"8b",x"c1",x"87"),
   870 => (x"c5",x"c8",x"48",x"d0"),
   871 => (x"7c",x"d5",x"c1",x"78"),
   872 => (x"31",x"c6",x"49",x"73"),
   873 => (x"97",x"d0",x"de",x"c2"),
   874 => (x"71",x"48",x"4a",x"bf"),
   875 => (x"ff",x"7c",x"70",x"b0"),
   876 => (x"78",x"c4",x"48",x"d0"),
   877 => (x"d5",x"fe",x"48",x"73"),
   878 => (x"5b",x"5e",x"0e",x"87"),
   879 => (x"f8",x"0e",x"5d",x"5c"),
   880 => (x"c0",x"4c",x"71",x"86"),
   881 => (x"87",x"e4",x"fb",x"7e"),
   882 => (x"f9",x"c0",x"4b",x"c0"),
   883 => (x"49",x"bf",x"97",x"e6"),
   884 => (x"cf",x"04",x"a9",x"c0"),
   885 => (x"87",x"f9",x"fb",x"87"),
   886 => (x"f9",x"c0",x"83",x"c1"),
   887 => (x"49",x"bf",x"97",x"e6"),
   888 => (x"87",x"f1",x"06",x"ab"),
   889 => (x"97",x"e6",x"f9",x"c0"),
   890 => (x"87",x"cf",x"02",x"bf"),
   891 => (x"70",x"87",x"f2",x"fa"),
   892 => (x"c6",x"02",x"99",x"49"),
   893 => (x"a9",x"ec",x"c0",x"87"),
   894 => (x"c0",x"87",x"f1",x"05"),
   895 => (x"87",x"e1",x"fa",x"4b"),
   896 => (x"dc",x"fa",x"4d",x"70"),
   897 => (x"58",x"a6",x"c8",x"87"),
   898 => (x"70",x"87",x"d6",x"fa"),
   899 => (x"c8",x"83",x"c1",x"4a"),
   900 => (x"69",x"97",x"49",x"a4"),
   901 => (x"c7",x"02",x"ad",x"49"),
   902 => (x"ad",x"ff",x"c0",x"87"),
   903 => (x"87",x"e7",x"c0",x"05"),
   904 => (x"97",x"49",x"a4",x"c9"),
   905 => (x"66",x"c4",x"49",x"69"),
   906 => (x"87",x"c7",x"02",x"a9"),
   907 => (x"a8",x"ff",x"c0",x"48"),
   908 => (x"ca",x"87",x"d4",x"05"),
   909 => (x"69",x"97",x"49",x"a4"),
   910 => (x"c6",x"02",x"aa",x"49"),
   911 => (x"aa",x"ff",x"c0",x"87"),
   912 => (x"c1",x"87",x"c4",x"05"),
   913 => (x"c0",x"87",x"d0",x"7e"),
   914 => (x"c6",x"02",x"ad",x"ec"),
   915 => (x"ad",x"fb",x"c0",x"87"),
   916 => (x"c0",x"87",x"c4",x"05"),
   917 => (x"6e",x"7e",x"c1",x"4b"),
   918 => (x"87",x"e1",x"fe",x"02"),
   919 => (x"73",x"87",x"e9",x"f9"),
   920 => (x"fb",x"8e",x"f8",x"48"),
   921 => (x"0e",x"00",x"87",x"e6"),
   922 => (x"5d",x"5c",x"5b",x"5e"),
   923 => (x"4b",x"71",x"1e",x"0e"),
   924 => (x"ab",x"4d",x"4c",x"c0"),
   925 => (x"87",x"e8",x"c0",x"04"),
   926 => (x"1e",x"f9",x"f6",x"c0"),
   927 => (x"c4",x"02",x"9d",x"75"),
   928 => (x"c2",x"4a",x"c0",x"87"),
   929 => (x"72",x"4a",x"c1",x"87"),
   930 => (x"87",x"e0",x"f0",x"49"),
   931 => (x"7e",x"70",x"86",x"c4"),
   932 => (x"05",x"6e",x"84",x"c1"),
   933 => (x"4c",x"73",x"87",x"c2"),
   934 => (x"ac",x"73",x"85",x"c1"),
   935 => (x"87",x"d8",x"ff",x"06"),
   936 => (x"26",x"26",x"48",x"6e"),
   937 => (x"26",x"4c",x"26",x"4d"),
   938 => (x"0e",x"4f",x"26",x"4b"),
   939 => (x"5d",x"5c",x"5b",x"5e"),
   940 => (x"4c",x"71",x"1e",x"0e"),
   941 => (x"c2",x"91",x"de",x"49"),
   942 => (x"71",x"4d",x"f1",x"ec"),
   943 => (x"02",x"6d",x"97",x"85"),
   944 => (x"c2",x"87",x"dd",x"c1"),
   945 => (x"4a",x"bf",x"dc",x"ec"),
   946 => (x"49",x"72",x"82",x"74"),
   947 => (x"70",x"87",x"d8",x"fe"),
   948 => (x"c0",x"02",x"6e",x"7e"),
   949 => (x"ec",x"c2",x"87",x"f3"),
   950 => (x"4a",x"6e",x"4b",x"e4"),
   951 => (x"c7",x"ff",x"49",x"cb"),
   952 => (x"4b",x"74",x"87",x"c6"),
   953 => (x"dd",x"c1",x"93",x"cb"),
   954 => (x"83",x"c4",x"83",x"fc"),
   955 => (x"7b",x"e4",x"fc",x"c0"),
   956 => (x"c3",x"c1",x"49",x"74"),
   957 => (x"7b",x"75",x"87",x"f5"),
   958 => (x"97",x"f0",x"ec",x"c2"),
   959 => (x"c2",x"1e",x"49",x"bf"),
   960 => (x"c1",x"49",x"e4",x"ec"),
   961 => (x"c4",x"87",x"cb",x"e1"),
   962 => (x"c1",x"49",x"74",x"86"),
   963 => (x"c0",x"87",x"dc",x"c3"),
   964 => (x"fb",x"c4",x"c1",x"49"),
   965 => (x"d8",x"ec",x"c2",x"87"),
   966 => (x"c1",x"78",x"c0",x"48"),
   967 => (x"87",x"d1",x"dd",x"49"),
   968 => (x"87",x"ff",x"fd",x"26"),
   969 => (x"64",x"61",x"6f",x"4c"),
   970 => (x"2e",x"67",x"6e",x"69"),
   971 => (x"0e",x"00",x"2e",x"2e"),
   972 => (x"0e",x"5c",x"5b",x"5e"),
   973 => (x"c2",x"4a",x"4b",x"71"),
   974 => (x"82",x"bf",x"dc",x"ec"),
   975 => (x"e6",x"fc",x"49",x"72"),
   976 => (x"9c",x"4c",x"70",x"87"),
   977 => (x"49",x"87",x"c4",x"02"),
   978 => (x"c2",x"87",x"e9",x"ec"),
   979 => (x"c0",x"48",x"dc",x"ec"),
   980 => (x"dc",x"49",x"c1",x"78"),
   981 => (x"cc",x"fd",x"87",x"db"),
   982 => (x"5b",x"5e",x"0e",x"87"),
   983 => (x"f4",x"0e",x"5d",x"5c"),
   984 => (x"e6",x"df",x"c2",x"86"),
   985 => (x"c4",x"4c",x"c0",x"4d"),
   986 => (x"78",x"c0",x"48",x"a6"),
   987 => (x"bf",x"dc",x"ec",x"c2"),
   988 => (x"06",x"a9",x"c0",x"49"),
   989 => (x"c2",x"87",x"c1",x"c1"),
   990 => (x"98",x"48",x"e6",x"df"),
   991 => (x"87",x"f8",x"c0",x"02"),
   992 => (x"1e",x"f9",x"f6",x"c0"),
   993 => (x"c7",x"02",x"66",x"c8"),
   994 => (x"48",x"a6",x"c4",x"87"),
   995 => (x"87",x"c5",x"78",x"c0"),
   996 => (x"c1",x"48",x"a6",x"c4"),
   997 => (x"49",x"66",x"c4",x"78"),
   998 => (x"c4",x"87",x"d1",x"ec"),
   999 => (x"c1",x"4d",x"70",x"86"),
  1000 => (x"48",x"66",x"c4",x"84"),
  1001 => (x"a6",x"c8",x"80",x"c1"),
  1002 => (x"dc",x"ec",x"c2",x"58"),
  1003 => (x"03",x"ac",x"49",x"bf"),
  1004 => (x"9d",x"75",x"87",x"c6"),
  1005 => (x"87",x"c8",x"ff",x"05"),
  1006 => (x"9d",x"75",x"4c",x"c0"),
  1007 => (x"87",x"e0",x"c3",x"02"),
  1008 => (x"1e",x"f9",x"f6",x"c0"),
  1009 => (x"c7",x"02",x"66",x"c8"),
  1010 => (x"48",x"a6",x"cc",x"87"),
  1011 => (x"87",x"c5",x"78",x"c0"),
  1012 => (x"c1",x"48",x"a6",x"cc"),
  1013 => (x"49",x"66",x"cc",x"78"),
  1014 => (x"c4",x"87",x"d1",x"eb"),
  1015 => (x"6e",x"7e",x"70",x"86"),
  1016 => (x"87",x"e9",x"c2",x"02"),
  1017 => (x"81",x"cb",x"49",x"6e"),
  1018 => (x"d0",x"49",x"69",x"97"),
  1019 => (x"d6",x"c1",x"02",x"99"),
  1020 => (x"ef",x"fc",x"c0",x"87"),
  1021 => (x"cb",x"49",x"74",x"4a"),
  1022 => (x"fc",x"dd",x"c1",x"91"),
  1023 => (x"c8",x"79",x"72",x"81"),
  1024 => (x"51",x"ff",x"c3",x"81"),
  1025 => (x"91",x"de",x"49",x"74"),
  1026 => (x"4d",x"f1",x"ec",x"c2"),
  1027 => (x"c1",x"c2",x"85",x"71"),
  1028 => (x"a5",x"c1",x"7d",x"97"),
  1029 => (x"51",x"e0",x"c0",x"49"),
  1030 => (x"97",x"f6",x"e7",x"c2"),
  1031 => (x"87",x"d2",x"02",x"bf"),
  1032 => (x"a5",x"c2",x"84",x"c1"),
  1033 => (x"f6",x"e7",x"c2",x"4b"),
  1034 => (x"ff",x"49",x"db",x"4a"),
  1035 => (x"c1",x"87",x"f9",x"c1"),
  1036 => (x"a5",x"cd",x"87",x"db"),
  1037 => (x"c1",x"51",x"c0",x"49"),
  1038 => (x"4b",x"a5",x"c2",x"84"),
  1039 => (x"49",x"cb",x"4a",x"6e"),
  1040 => (x"87",x"e4",x"c1",x"ff"),
  1041 => (x"c0",x"87",x"c6",x"c1"),
  1042 => (x"74",x"4a",x"eb",x"fa"),
  1043 => (x"c1",x"91",x"cb",x"49"),
  1044 => (x"72",x"81",x"fc",x"dd"),
  1045 => (x"f6",x"e7",x"c2",x"79"),
  1046 => (x"d8",x"02",x"bf",x"97"),
  1047 => (x"de",x"49",x"74",x"87"),
  1048 => (x"c2",x"84",x"c1",x"91"),
  1049 => (x"71",x"4b",x"f1",x"ec"),
  1050 => (x"f6",x"e7",x"c2",x"83"),
  1051 => (x"ff",x"49",x"dd",x"4a"),
  1052 => (x"d8",x"87",x"f5",x"c0"),
  1053 => (x"de",x"4b",x"74",x"87"),
  1054 => (x"f1",x"ec",x"c2",x"93"),
  1055 => (x"49",x"a3",x"cb",x"83"),
  1056 => (x"84",x"c1",x"51",x"c0"),
  1057 => (x"cb",x"4a",x"6e",x"73"),
  1058 => (x"db",x"c0",x"ff",x"49"),
  1059 => (x"48",x"66",x"c4",x"87"),
  1060 => (x"a6",x"c8",x"80",x"c1"),
  1061 => (x"03",x"ac",x"c7",x"58"),
  1062 => (x"6e",x"87",x"c5",x"c0"),
  1063 => (x"87",x"e0",x"fc",x"05"),
  1064 => (x"8e",x"f4",x"48",x"74"),
  1065 => (x"1e",x"87",x"fc",x"f7"),
  1066 => (x"4b",x"71",x"1e",x"73"),
  1067 => (x"c1",x"91",x"cb",x"49"),
  1068 => (x"c8",x"81",x"fc",x"dd"),
  1069 => (x"de",x"c2",x"4a",x"a1"),
  1070 => (x"50",x"12",x"48",x"d0"),
  1071 => (x"c0",x"4a",x"a1",x"c9"),
  1072 => (x"12",x"48",x"e6",x"f9"),
  1073 => (x"c2",x"81",x"ca",x"50"),
  1074 => (x"11",x"48",x"f0",x"ec"),
  1075 => (x"f0",x"ec",x"c2",x"50"),
  1076 => (x"1e",x"49",x"bf",x"97"),
  1077 => (x"d9",x"c1",x"49",x"c0"),
  1078 => (x"ec",x"c2",x"87",x"f8"),
  1079 => (x"78",x"de",x"48",x"d8"),
  1080 => (x"cc",x"d6",x"49",x"c1"),
  1081 => (x"fe",x"f6",x"26",x"87"),
  1082 => (x"4a",x"71",x"1e",x"87"),
  1083 => (x"c1",x"91",x"cb",x"49"),
  1084 => (x"c8",x"81",x"fc",x"dd"),
  1085 => (x"c2",x"48",x"11",x"81"),
  1086 => (x"c2",x"58",x"dc",x"ec"),
  1087 => (x"c0",x"48",x"dc",x"ec"),
  1088 => (x"d5",x"49",x"c1",x"78"),
  1089 => (x"4f",x"26",x"87",x"eb"),
  1090 => (x"c0",x"49",x"c0",x"1e"),
  1091 => (x"26",x"87",x"c1",x"fd"),
  1092 => (x"99",x"71",x"1e",x"4f"),
  1093 => (x"c1",x"87",x"d2",x"02"),
  1094 => (x"c0",x"48",x"d1",x"df"),
  1095 => (x"c1",x"80",x"f7",x"50"),
  1096 => (x"c1",x"40",x"e9",x"c3"),
  1097 => (x"ce",x"78",x"f5",x"dd"),
  1098 => (x"cd",x"df",x"c1",x"87"),
  1099 => (x"ee",x"dd",x"c1",x"48"),
  1100 => (x"c1",x"80",x"fc",x"78"),
  1101 => (x"26",x"78",x"c8",x"c4"),
  1102 => (x"5b",x"5e",x"0e",x"4f"),
  1103 => (x"4c",x"71",x"0e",x"5c"),
  1104 => (x"c1",x"92",x"cb",x"4a"),
  1105 => (x"c8",x"82",x"fc",x"dd"),
  1106 => (x"a2",x"c9",x"49",x"a2"),
  1107 => (x"4b",x"6b",x"97",x"4b"),
  1108 => (x"49",x"69",x"97",x"1e"),
  1109 => (x"12",x"82",x"ca",x"1e"),
  1110 => (x"fc",x"e7",x"c0",x"49"),
  1111 => (x"d4",x"49",x"c0",x"87"),
  1112 => (x"49",x"74",x"87",x"cf"),
  1113 => (x"87",x"c3",x"fa",x"c0"),
  1114 => (x"f8",x"f4",x"8e",x"f8"),
  1115 => (x"1e",x"73",x"1e",x"87"),
  1116 => (x"ff",x"49",x"4b",x"71"),
  1117 => (x"49",x"73",x"87",x"c3"),
  1118 => (x"c0",x"87",x"fe",x"fe"),
  1119 => (x"cf",x"fb",x"c0",x"49"),
  1120 => (x"87",x"e3",x"f4",x"87"),
  1121 => (x"71",x"1e",x"73",x"1e"),
  1122 => (x"4a",x"a3",x"c6",x"4b"),
  1123 => (x"c1",x"87",x"db",x"02"),
  1124 => (x"87",x"d6",x"02",x"8a"),
  1125 => (x"da",x"c1",x"02",x"8a"),
  1126 => (x"c0",x"02",x"8a",x"87"),
  1127 => (x"02",x"8a",x"87",x"fc"),
  1128 => (x"8a",x"87",x"e1",x"c0"),
  1129 => (x"c1",x"87",x"cb",x"02"),
  1130 => (x"49",x"c7",x"87",x"db"),
  1131 => (x"c1",x"87",x"fa",x"fc"),
  1132 => (x"ec",x"c2",x"87",x"de"),
  1133 => (x"c1",x"02",x"bf",x"dc"),
  1134 => (x"c1",x"48",x"87",x"cb"),
  1135 => (x"e0",x"ec",x"c2",x"88"),
  1136 => (x"87",x"c1",x"c1",x"58"),
  1137 => (x"bf",x"e0",x"ec",x"c2"),
  1138 => (x"87",x"f9",x"c0",x"02"),
  1139 => (x"bf",x"dc",x"ec",x"c2"),
  1140 => (x"c2",x"80",x"c1",x"48"),
  1141 => (x"c0",x"58",x"e0",x"ec"),
  1142 => (x"ec",x"c2",x"87",x"eb"),
  1143 => (x"c6",x"49",x"bf",x"dc"),
  1144 => (x"e0",x"ec",x"c2",x"89"),
  1145 => (x"a9",x"b7",x"c0",x"59"),
  1146 => (x"c2",x"87",x"da",x"03"),
  1147 => (x"c0",x"48",x"dc",x"ec"),
  1148 => (x"c2",x"87",x"d2",x"78"),
  1149 => (x"02",x"bf",x"e0",x"ec"),
  1150 => (x"ec",x"c2",x"87",x"cb"),
  1151 => (x"c6",x"48",x"bf",x"dc"),
  1152 => (x"e0",x"ec",x"c2",x"80"),
  1153 => (x"d1",x"49",x"c0",x"58"),
  1154 => (x"49",x"73",x"87",x"e7"),
  1155 => (x"87",x"db",x"f7",x"c0"),
  1156 => (x"0e",x"87",x"d4",x"f2"),
  1157 => (x"0e",x"5c",x"5b",x"5e"),
  1158 => (x"66",x"cc",x"4c",x"71"),
  1159 => (x"cb",x"4b",x"74",x"1e"),
  1160 => (x"fc",x"dd",x"c1",x"93"),
  1161 => (x"4a",x"a3",x"c4",x"83"),
  1162 => (x"fa",x"fe",x"49",x"6a"),
  1163 => (x"c2",x"c1",x"87",x"ca"),
  1164 => (x"a3",x"c8",x"7b",x"e7"),
  1165 => (x"51",x"66",x"d4",x"49"),
  1166 => (x"d8",x"49",x"a3",x"c9"),
  1167 => (x"a3",x"ca",x"51",x"66"),
  1168 => (x"51",x"66",x"dc",x"49"),
  1169 => (x"87",x"dd",x"f1",x"26"),
  1170 => (x"5c",x"5b",x"5e",x"0e"),
  1171 => (x"d0",x"ff",x"0e",x"5d"),
  1172 => (x"59",x"a6",x"d8",x"86"),
  1173 => (x"c0",x"48",x"a6",x"c4"),
  1174 => (x"c1",x"80",x"c4",x"78"),
  1175 => (x"c4",x"78",x"66",x"c4"),
  1176 => (x"c4",x"78",x"c1",x"80"),
  1177 => (x"c2",x"78",x"c1",x"80"),
  1178 => (x"c1",x"48",x"e0",x"ec"),
  1179 => (x"d8",x"ec",x"c2",x"78"),
  1180 => (x"a8",x"de",x"48",x"bf"),
  1181 => (x"f3",x"87",x"cb",x"05"),
  1182 => (x"49",x"70",x"87",x"df"),
  1183 => (x"ce",x"59",x"a6",x"c8"),
  1184 => (x"e7",x"e8",x"87",x"f8"),
  1185 => (x"87",x"c9",x"e9",x"87"),
  1186 => (x"70",x"87",x"d6",x"e8"),
  1187 => (x"ac",x"fb",x"c0",x"4c"),
  1188 => (x"87",x"d0",x"c1",x"02"),
  1189 => (x"c1",x"05",x"66",x"d4"),
  1190 => (x"1e",x"c0",x"87",x"c2"),
  1191 => (x"c1",x"1e",x"c1",x"1e"),
  1192 => (x"c0",x"1e",x"ef",x"df"),
  1193 => (x"87",x"eb",x"fd",x"49"),
  1194 => (x"4a",x"66",x"d0",x"c1"),
  1195 => (x"49",x"6a",x"82",x"c4"),
  1196 => (x"51",x"74",x"81",x"c7"),
  1197 => (x"1e",x"d8",x"1e",x"c1"),
  1198 => (x"81",x"c8",x"49",x"6a"),
  1199 => (x"d8",x"87",x"e6",x"e8"),
  1200 => (x"66",x"c4",x"c1",x"86"),
  1201 => (x"01",x"a8",x"c0",x"48"),
  1202 => (x"a6",x"c4",x"87",x"c7"),
  1203 => (x"ce",x"78",x"c1",x"48"),
  1204 => (x"66",x"c4",x"c1",x"87"),
  1205 => (x"cc",x"88",x"c1",x"48"),
  1206 => (x"87",x"c3",x"58",x"a6"),
  1207 => (x"cc",x"87",x"f2",x"e7"),
  1208 => (x"78",x"c2",x"48",x"a6"),
  1209 => (x"cd",x"02",x"9c",x"74"),
  1210 => (x"66",x"c4",x"87",x"cc"),
  1211 => (x"66",x"c8",x"c1",x"48"),
  1212 => (x"c1",x"cd",x"03",x"a8"),
  1213 => (x"48",x"a6",x"d8",x"87"),
  1214 => (x"e4",x"e6",x"78",x"c0"),
  1215 => (x"c1",x"4c",x"70",x"87"),
  1216 => (x"c2",x"05",x"ac",x"d0"),
  1217 => (x"66",x"d8",x"87",x"d6"),
  1218 => (x"87",x"c8",x"e9",x"7e"),
  1219 => (x"a6",x"dc",x"49",x"70"),
  1220 => (x"87",x"cd",x"e6",x"59"),
  1221 => (x"ec",x"c0",x"4c",x"70"),
  1222 => (x"ea",x"c1",x"05",x"ac"),
  1223 => (x"49",x"66",x"c4",x"87"),
  1224 => (x"c0",x"c1",x"91",x"cb"),
  1225 => (x"a1",x"c4",x"81",x"66"),
  1226 => (x"c8",x"4d",x"6a",x"4a"),
  1227 => (x"66",x"d8",x"4a",x"a1"),
  1228 => (x"e9",x"c3",x"c1",x"52"),
  1229 => (x"87",x"e9",x"e5",x"79"),
  1230 => (x"02",x"9c",x"4c",x"70"),
  1231 => (x"fb",x"c0",x"87",x"d8"),
  1232 => (x"87",x"d2",x"02",x"ac"),
  1233 => (x"d8",x"e5",x"55",x"74"),
  1234 => (x"9c",x"4c",x"70",x"87"),
  1235 => (x"c0",x"87",x"c7",x"02"),
  1236 => (x"ff",x"05",x"ac",x"fb"),
  1237 => (x"e0",x"c0",x"87",x"ee"),
  1238 => (x"55",x"c1",x"c2",x"55"),
  1239 => (x"d4",x"7d",x"97",x"c0"),
  1240 => (x"a9",x"6e",x"49",x"66"),
  1241 => (x"c4",x"87",x"db",x"05"),
  1242 => (x"66",x"c8",x"48",x"66"),
  1243 => (x"87",x"ca",x"04",x"a8"),
  1244 => (x"c1",x"48",x"66",x"c4"),
  1245 => (x"58",x"a6",x"c8",x"80"),
  1246 => (x"66",x"c8",x"87",x"c8"),
  1247 => (x"cc",x"88",x"c1",x"48"),
  1248 => (x"dc",x"e4",x"58",x"a6"),
  1249 => (x"c1",x"4c",x"70",x"87"),
  1250 => (x"c8",x"05",x"ac",x"d0"),
  1251 => (x"48",x"66",x"d0",x"87"),
  1252 => (x"a6",x"d4",x"80",x"c1"),
  1253 => (x"ac",x"d0",x"c1",x"58"),
  1254 => (x"87",x"ea",x"fd",x"02"),
  1255 => (x"d4",x"48",x"a6",x"dc"),
  1256 => (x"66",x"d8",x"78",x"66"),
  1257 => (x"a8",x"66",x"dc",x"48"),
  1258 => (x"87",x"dc",x"c9",x"05"),
  1259 => (x"48",x"a6",x"e0",x"c0"),
  1260 => (x"c4",x"78",x"f0",x"c0"),
  1261 => (x"78",x"66",x"cc",x"80"),
  1262 => (x"78",x"c0",x"80",x"c4"),
  1263 => (x"c0",x"48",x"74",x"7e"),
  1264 => (x"f0",x"c0",x"88",x"fb"),
  1265 => (x"98",x"70",x"58",x"a6"),
  1266 => (x"87",x"d7",x"c8",x"02"),
  1267 => (x"c0",x"88",x"cb",x"48"),
  1268 => (x"70",x"58",x"a6",x"f0"),
  1269 => (x"e9",x"c0",x"02",x"98"),
  1270 => (x"88",x"c9",x"48",x"87"),
  1271 => (x"58",x"a6",x"f0",x"c0"),
  1272 => (x"c3",x"02",x"98",x"70"),
  1273 => (x"c4",x"48",x"87",x"e1"),
  1274 => (x"a6",x"f0",x"c0",x"88"),
  1275 => (x"02",x"98",x"70",x"58"),
  1276 => (x"c1",x"48",x"87",x"de"),
  1277 => (x"a6",x"f0",x"c0",x"88"),
  1278 => (x"02",x"98",x"70",x"58"),
  1279 => (x"c7",x"87",x"c8",x"c3"),
  1280 => (x"e0",x"c0",x"87",x"db"),
  1281 => (x"78",x"c0",x"48",x"a6"),
  1282 => (x"c1",x"48",x"66",x"cc"),
  1283 => (x"58",x"a6",x"d0",x"80"),
  1284 => (x"70",x"87",x"ce",x"e2"),
  1285 => (x"ac",x"ec",x"c0",x"4c"),
  1286 => (x"c0",x"87",x"d5",x"02"),
  1287 => (x"c6",x"02",x"66",x"e0"),
  1288 => (x"a6",x"e4",x"c0",x"87"),
  1289 => (x"74",x"87",x"c9",x"5c"),
  1290 => (x"88",x"f0",x"c0",x"48"),
  1291 => (x"58",x"a6",x"e8",x"c0"),
  1292 => (x"02",x"ac",x"ec",x"c0"),
  1293 => (x"e8",x"e1",x"87",x"cc"),
  1294 => (x"c0",x"4c",x"70",x"87"),
  1295 => (x"ff",x"05",x"ac",x"ec"),
  1296 => (x"e0",x"c0",x"87",x"f4"),
  1297 => (x"66",x"d4",x"1e",x"66"),
  1298 => (x"ec",x"c0",x"1e",x"49"),
  1299 => (x"df",x"c1",x"1e",x"66"),
  1300 => (x"66",x"d4",x"1e",x"ef"),
  1301 => (x"87",x"fb",x"f6",x"49"),
  1302 => (x"1e",x"ca",x"1e",x"c0"),
  1303 => (x"cb",x"49",x"66",x"dc"),
  1304 => (x"66",x"d8",x"c1",x"91"),
  1305 => (x"48",x"a6",x"d8",x"81"),
  1306 => (x"d8",x"78",x"a1",x"c4"),
  1307 => (x"e1",x"49",x"bf",x"66"),
  1308 => (x"86",x"d8",x"87",x"f3"),
  1309 => (x"06",x"a8",x"b7",x"c0"),
  1310 => (x"c1",x"87",x"c7",x"c1"),
  1311 => (x"c8",x"1e",x"de",x"1e"),
  1312 => (x"e1",x"49",x"bf",x"66"),
  1313 => (x"86",x"c8",x"87",x"df"),
  1314 => (x"c0",x"48",x"49",x"70"),
  1315 => (x"e4",x"c0",x"88",x"08"),
  1316 => (x"b7",x"c0",x"58",x"a6"),
  1317 => (x"e9",x"c0",x"06",x"a8"),
  1318 => (x"66",x"e0",x"c0",x"87"),
  1319 => (x"a8",x"b7",x"dd",x"48"),
  1320 => (x"6e",x"87",x"df",x"03"),
  1321 => (x"e0",x"c0",x"49",x"bf"),
  1322 => (x"e0",x"c0",x"81",x"66"),
  1323 => (x"c1",x"49",x"66",x"51"),
  1324 => (x"81",x"bf",x"6e",x"81"),
  1325 => (x"c0",x"51",x"c1",x"c2"),
  1326 => (x"c2",x"49",x"66",x"e0"),
  1327 => (x"81",x"bf",x"6e",x"81"),
  1328 => (x"7e",x"c1",x"51",x"c0"),
  1329 => (x"e2",x"87",x"dc",x"c4"),
  1330 => (x"e4",x"c0",x"87",x"ca"),
  1331 => (x"c3",x"e2",x"58",x"a6"),
  1332 => (x"a6",x"e8",x"c0",x"87"),
  1333 => (x"a8",x"ec",x"c0",x"58"),
  1334 => (x"87",x"cb",x"c0",x"05"),
  1335 => (x"48",x"a6",x"e4",x"c0"),
  1336 => (x"78",x"66",x"e0",x"c0"),
  1337 => (x"ff",x"87",x"c4",x"c0"),
  1338 => (x"c4",x"87",x"f6",x"de"),
  1339 => (x"91",x"cb",x"49",x"66"),
  1340 => (x"48",x"66",x"c0",x"c1"),
  1341 => (x"7e",x"70",x"80",x"71"),
  1342 => (x"82",x"c8",x"4a",x"6e"),
  1343 => (x"81",x"ca",x"49",x"6e"),
  1344 => (x"51",x"66",x"e0",x"c0"),
  1345 => (x"49",x"66",x"e4",x"c0"),
  1346 => (x"e0",x"c0",x"81",x"c1"),
  1347 => (x"48",x"c1",x"89",x"66"),
  1348 => (x"49",x"70",x"30",x"71"),
  1349 => (x"97",x"71",x"89",x"c1"),
  1350 => (x"cd",x"f0",x"c2",x"7a"),
  1351 => (x"e0",x"c0",x"49",x"bf"),
  1352 => (x"6a",x"97",x"29",x"66"),
  1353 => (x"98",x"71",x"48",x"4a"),
  1354 => (x"58",x"a6",x"f0",x"c0"),
  1355 => (x"81",x"c4",x"49",x"6e"),
  1356 => (x"66",x"dc",x"4d",x"69"),
  1357 => (x"a8",x"66",x"d8",x"48"),
  1358 => (x"87",x"c8",x"c0",x"02"),
  1359 => (x"c0",x"48",x"a6",x"d8"),
  1360 => (x"87",x"c5",x"c0",x"78"),
  1361 => (x"c1",x"48",x"a6",x"d8"),
  1362 => (x"1e",x"66",x"d8",x"78"),
  1363 => (x"75",x"1e",x"e0",x"c0"),
  1364 => (x"d0",x"de",x"ff",x"49"),
  1365 => (x"70",x"86",x"c8",x"87"),
  1366 => (x"ac",x"b7",x"c0",x"4c"),
  1367 => (x"87",x"d4",x"c1",x"06"),
  1368 => (x"e0",x"c0",x"85",x"74"),
  1369 => (x"75",x"89",x"74",x"49"),
  1370 => (x"ee",x"d9",x"c1",x"4b"),
  1371 => (x"ec",x"fe",x"71",x"4a"),
  1372 => (x"85",x"c2",x"87",x"f6"),
  1373 => (x"48",x"66",x"e8",x"c0"),
  1374 => (x"ec",x"c0",x"80",x"c1"),
  1375 => (x"ec",x"c0",x"58",x"a6"),
  1376 => (x"81",x"c1",x"49",x"66"),
  1377 => (x"c0",x"02",x"a9",x"70"),
  1378 => (x"a6",x"d8",x"87",x"c8"),
  1379 => (x"c0",x"78",x"c0",x"48"),
  1380 => (x"a6",x"d8",x"87",x"c5"),
  1381 => (x"d8",x"78",x"c1",x"48"),
  1382 => (x"a4",x"c2",x"1e",x"66"),
  1383 => (x"48",x"e0",x"c0",x"49"),
  1384 => (x"49",x"70",x"88",x"71"),
  1385 => (x"ff",x"49",x"75",x"1e"),
  1386 => (x"c8",x"87",x"fa",x"dc"),
  1387 => (x"a8",x"b7",x"c0",x"86"),
  1388 => (x"87",x"c0",x"ff",x"01"),
  1389 => (x"02",x"66",x"e8",x"c0"),
  1390 => (x"6e",x"87",x"d1",x"c0"),
  1391 => (x"c0",x"81",x"c9",x"49"),
  1392 => (x"6e",x"51",x"66",x"e8"),
  1393 => (x"f9",x"c4",x"c1",x"48"),
  1394 => (x"87",x"cc",x"c0",x"78"),
  1395 => (x"81",x"c9",x"49",x"6e"),
  1396 => (x"48",x"6e",x"51",x"c2"),
  1397 => (x"78",x"ed",x"c5",x"c1"),
  1398 => (x"c6",x"c0",x"7e",x"c1"),
  1399 => (x"f0",x"db",x"ff",x"87"),
  1400 => (x"6e",x"4c",x"70",x"87"),
  1401 => (x"87",x"f5",x"c0",x"02"),
  1402 => (x"c8",x"48",x"66",x"c4"),
  1403 => (x"c0",x"04",x"a8",x"66"),
  1404 => (x"66",x"c4",x"87",x"cb"),
  1405 => (x"c8",x"80",x"c1",x"48"),
  1406 => (x"e0",x"c0",x"58",x"a6"),
  1407 => (x"48",x"66",x"c8",x"87"),
  1408 => (x"a6",x"cc",x"88",x"c1"),
  1409 => (x"87",x"d5",x"c0",x"58"),
  1410 => (x"05",x"ac",x"c6",x"c1"),
  1411 => (x"cc",x"87",x"c8",x"c0"),
  1412 => (x"80",x"c1",x"48",x"66"),
  1413 => (x"ff",x"58",x"a6",x"d0"),
  1414 => (x"70",x"87",x"f6",x"da"),
  1415 => (x"48",x"66",x"d0",x"4c"),
  1416 => (x"a6",x"d4",x"80",x"c1"),
  1417 => (x"02",x"9c",x"74",x"58"),
  1418 => (x"c4",x"87",x"cb",x"c0"),
  1419 => (x"c8",x"c1",x"48",x"66"),
  1420 => (x"f2",x"04",x"a8",x"66"),
  1421 => (x"da",x"ff",x"87",x"ff"),
  1422 => (x"66",x"c4",x"87",x"ce"),
  1423 => (x"03",x"a8",x"c7",x"48"),
  1424 => (x"c2",x"87",x"e5",x"c0"),
  1425 => (x"c0",x"48",x"e0",x"ec"),
  1426 => (x"49",x"66",x"c4",x"78"),
  1427 => (x"c0",x"c1",x"91",x"cb"),
  1428 => (x"a1",x"c4",x"81",x"66"),
  1429 => (x"c0",x"4a",x"6a",x"4a"),
  1430 => (x"66",x"c4",x"79",x"52"),
  1431 => (x"c8",x"80",x"c1",x"48"),
  1432 => (x"a8",x"c7",x"58",x"a6"),
  1433 => (x"87",x"db",x"ff",x"04"),
  1434 => (x"e0",x"8e",x"d0",x"ff"),
  1435 => (x"20",x"3a",x"87",x"f5"),
  1436 => (x"1e",x"73",x"1e",x"00"),
  1437 => (x"02",x"9b",x"4b",x"71"),
  1438 => (x"ec",x"c2",x"87",x"c6"),
  1439 => (x"78",x"c0",x"48",x"dc"),
  1440 => (x"ec",x"c2",x"1e",x"c7"),
  1441 => (x"1e",x"49",x"bf",x"dc"),
  1442 => (x"1e",x"fc",x"dd",x"c1"),
  1443 => (x"bf",x"d8",x"ec",x"c2"),
  1444 => (x"87",x"f4",x"ee",x"49"),
  1445 => (x"ec",x"c2",x"86",x"cc"),
  1446 => (x"e9",x"49",x"bf",x"d8"),
  1447 => (x"9b",x"73",x"87",x"f3"),
  1448 => (x"c1",x"87",x"c8",x"02"),
  1449 => (x"c0",x"49",x"fc",x"dd"),
  1450 => (x"ff",x"87",x"d2",x"e6"),
  1451 => (x"1e",x"87",x"f8",x"df"),
  1452 => (x"4b",x"c0",x"1e",x"73"),
  1453 => (x"48",x"d0",x"de",x"c2"),
  1454 => (x"df",x"c1",x"50",x"c0"),
  1455 => (x"c0",x"49",x"bf",x"df"),
  1456 => (x"70",x"87",x"e2",x"fe"),
  1457 => (x"87",x"c4",x"05",x"98"),
  1458 => (x"4b",x"d2",x"db",x"c1"),
  1459 => (x"df",x"ff",x"48",x"73"),
  1460 => (x"4f",x"52",x"87",x"d5"),
  1461 => (x"6f",x"6c",x"20",x"4d"),
  1462 => (x"6e",x"69",x"64",x"61"),
  1463 => (x"61",x"66",x"20",x"67"),
  1464 => (x"64",x"65",x"6c",x"69"),
  1465 => (x"e5",x"c7",x"1e",x"00"),
  1466 => (x"fe",x"49",x"c1",x"87"),
  1467 => (x"ef",x"fe",x"87",x"c3"),
  1468 => (x"98",x"70",x"87",x"c9"),
  1469 => (x"fe",x"87",x"cd",x"02"),
  1470 => (x"70",x"87",x"c6",x"f8"),
  1471 => (x"87",x"c4",x"02",x"98"),
  1472 => (x"87",x"c2",x"4a",x"c1"),
  1473 => (x"9a",x"72",x"4a",x"c0"),
  1474 => (x"c0",x"87",x"ce",x"05"),
  1475 => (x"f5",x"dc",x"c1",x"1e"),
  1476 => (x"de",x"f3",x"c0",x"49"),
  1477 => (x"fe",x"86",x"c4",x"87"),
  1478 => (x"c1",x"1e",x"c0",x"87"),
  1479 => (x"c0",x"49",x"c0",x"dd"),
  1480 => (x"c0",x"87",x"d0",x"f3"),
  1481 => (x"87",x"c7",x"fe",x"1e"),
  1482 => (x"f3",x"c0",x"49",x"70"),
  1483 => (x"dc",x"c3",x"87",x"c5"),
  1484 => (x"26",x"8e",x"f8",x"87"),
  1485 => (x"20",x"44",x"53",x"4f"),
  1486 => (x"6c",x"69",x"61",x"66"),
  1487 => (x"00",x"2e",x"64",x"65"),
  1488 => (x"74",x"6f",x"6f",x"42"),
  1489 => (x"2e",x"67",x"6e",x"69"),
  1490 => (x"1e",x"00",x"2e",x"2e"),
  1491 => (x"87",x"d0",x"e8",x"c0"),
  1492 => (x"87",x"ea",x"f6",x"c0"),
  1493 => (x"4f",x"26",x"87",x"f6"),
  1494 => (x"dc",x"ec",x"c2",x"1e"),
  1495 => (x"c2",x"78",x"c0",x"48"),
  1496 => (x"c0",x"48",x"d8",x"ec"),
  1497 => (x"87",x"fd",x"fd",x"78"),
  1498 => (x"48",x"c0",x"87",x"e1"),
  1499 => (x"20",x"80",x"4f",x"26"),
  1500 => (x"74",x"69",x"78",x"45"),
  1501 => (x"42",x"20",x"80",x"00"),
  1502 => (x"00",x"6b",x"63",x"61"),
  1503 => (x"00",x"00",x"10",x"e9"),
  1504 => (x"00",x"00",x"2b",x"31"),
  1505 => (x"e9",x"00",x"00",x"00"),
  1506 => (x"4f",x"00",x"00",x"10"),
  1507 => (x"00",x"00",x"00",x"2b"),
  1508 => (x"10",x"e9",x"00",x"00"),
  1509 => (x"2b",x"6d",x"00",x"00"),
  1510 => (x"00",x"00",x"00",x"00"),
  1511 => (x"00",x"10",x"e9",x"00"),
  1512 => (x"00",x"2b",x"8b",x"00"),
  1513 => (x"00",x"00",x"00",x"00"),
  1514 => (x"00",x"00",x"10",x"e9"),
  1515 => (x"00",x"00",x"2b",x"a9"),
  1516 => (x"e9",x"00",x"00",x"00"),
  1517 => (x"c7",x"00",x"00",x"10"),
  1518 => (x"00",x"00",x"00",x"2b"),
  1519 => (x"10",x"e9",x"00",x"00"),
  1520 => (x"2b",x"e5",x"00",x"00"),
  1521 => (x"00",x"00",x"00",x"00"),
  1522 => (x"00",x"10",x"e9",x"00"),
  1523 => (x"00",x"00",x"00",x"00"),
  1524 => (x"00",x"00",x"00",x"00"),
  1525 => (x"00",x"00",x"11",x"84"),
  1526 => (x"00",x"00",x"00",x"00"),
  1527 => (x"e3",x"00",x"00",x"00"),
  1528 => (x"43",x"00",x"00",x"17"),
  1529 => (x"20",x"20",x"36",x"31"),
  1530 => (x"52",x"20",x"20",x"20"),
  1531 => (x"4c",x"00",x"4d",x"4f"),
  1532 => (x"20",x"64",x"61",x"6f"),
  1533 => (x"1e",x"00",x"2e",x"2a"),
  1534 => (x"c0",x"48",x"f0",x"fe"),
  1535 => (x"79",x"09",x"cd",x"78"),
  1536 => (x"1e",x"4f",x"26",x"09"),
  1537 => (x"bf",x"f0",x"fe",x"1e"),
  1538 => (x"26",x"26",x"48",x"7e"),
  1539 => (x"f0",x"fe",x"1e",x"4f"),
  1540 => (x"26",x"78",x"c1",x"48"),
  1541 => (x"f0",x"fe",x"1e",x"4f"),
  1542 => (x"26",x"78",x"c0",x"48"),
  1543 => (x"4a",x"71",x"1e",x"4f"),
  1544 => (x"26",x"52",x"52",x"c0"),
  1545 => (x"5b",x"5e",x"0e",x"4f"),
  1546 => (x"f4",x"0e",x"5d",x"5c"),
  1547 => (x"97",x"4d",x"71",x"86"),
  1548 => (x"a5",x"c1",x"7e",x"6d"),
  1549 => (x"48",x"6c",x"97",x"4c"),
  1550 => (x"6e",x"58",x"a6",x"c8"),
  1551 => (x"a8",x"66",x"c4",x"48"),
  1552 => (x"ff",x"87",x"c5",x"05"),
  1553 => (x"87",x"e6",x"c0",x"48"),
  1554 => (x"c2",x"87",x"ca",x"ff"),
  1555 => (x"6c",x"97",x"49",x"a5"),
  1556 => (x"4b",x"a3",x"71",x"4b"),
  1557 => (x"97",x"4b",x"6b",x"97"),
  1558 => (x"48",x"6e",x"7e",x"6c"),
  1559 => (x"a6",x"c8",x"80",x"c1"),
  1560 => (x"cc",x"98",x"c7",x"58"),
  1561 => (x"97",x"70",x"58",x"a6"),
  1562 => (x"87",x"e1",x"fe",x"7c"),
  1563 => (x"8e",x"f4",x"48",x"73"),
  1564 => (x"4c",x"26",x"4d",x"26"),
  1565 => (x"4f",x"26",x"4b",x"26"),
  1566 => (x"5c",x"5b",x"5e",x"0e"),
  1567 => (x"71",x"86",x"f4",x"0e"),
  1568 => (x"4a",x"66",x"d8",x"4c"),
  1569 => (x"c2",x"9a",x"ff",x"c3"),
  1570 => (x"6c",x"97",x"4b",x"a4"),
  1571 => (x"49",x"a1",x"73",x"49"),
  1572 => (x"6c",x"97",x"51",x"72"),
  1573 => (x"c1",x"48",x"6e",x"7e"),
  1574 => (x"58",x"a6",x"c8",x"80"),
  1575 => (x"a6",x"cc",x"98",x"c7"),
  1576 => (x"f4",x"54",x"70",x"58"),
  1577 => (x"87",x"ca",x"ff",x"8e"),
  1578 => (x"e8",x"fd",x"1e",x"1e"),
  1579 => (x"4a",x"bf",x"e0",x"87"),
  1580 => (x"c0",x"e0",x"c0",x"49"),
  1581 => (x"87",x"cb",x"02",x"99"),
  1582 => (x"f0",x"c2",x"1e",x"72"),
  1583 => (x"f7",x"fe",x"49",x"c3"),
  1584 => (x"fc",x"86",x"c4",x"87"),
  1585 => (x"7e",x"70",x"87",x"fd"),
  1586 => (x"26",x"87",x"c2",x"fd"),
  1587 => (x"c2",x"1e",x"4f",x"26"),
  1588 => (x"fd",x"49",x"c3",x"f0"),
  1589 => (x"e2",x"c1",x"87",x"c7"),
  1590 => (x"da",x"fc",x"49",x"e8"),
  1591 => (x"87",x"d9",x"c5",x"87"),
  1592 => (x"5e",x"0e",x"4f",x"26"),
  1593 => (x"0e",x"5d",x"5c",x"5b"),
  1594 => (x"bf",x"e2",x"f0",x"c2"),
  1595 => (x"f6",x"e4",x"c1",x"4a"),
  1596 => (x"72",x"4c",x"49",x"bf"),
  1597 => (x"fc",x"4d",x"71",x"bc"),
  1598 => (x"4b",x"c0",x"87",x"db"),
  1599 => (x"99",x"d0",x"49",x"74"),
  1600 => (x"75",x"87",x"d5",x"02"),
  1601 => (x"71",x"99",x"d0",x"49"),
  1602 => (x"c1",x"1e",x"c0",x"1e"),
  1603 => (x"73",x"4a",x"c8",x"eb"),
  1604 => (x"c0",x"49",x"12",x"82"),
  1605 => (x"86",x"c8",x"87",x"e4"),
  1606 => (x"83",x"2d",x"2c",x"c1"),
  1607 => (x"ff",x"04",x"ab",x"c8"),
  1608 => (x"e8",x"fb",x"87",x"da"),
  1609 => (x"f6",x"e4",x"c1",x"87"),
  1610 => (x"e2",x"f0",x"c2",x"48"),
  1611 => (x"4d",x"26",x"78",x"bf"),
  1612 => (x"4b",x"26",x"4c",x"26"),
  1613 => (x"00",x"00",x"4f",x"26"),
  1614 => (x"ff",x"1e",x"00",x"00"),
  1615 => (x"e1",x"c8",x"48",x"d0"),
  1616 => (x"48",x"d4",x"ff",x"78"),
  1617 => (x"66",x"c4",x"78",x"c5"),
  1618 => (x"c3",x"87",x"c3",x"02"),
  1619 => (x"66",x"c8",x"78",x"e0"),
  1620 => (x"ff",x"87",x"c6",x"02"),
  1621 => (x"f0",x"c3",x"48",x"d4"),
  1622 => (x"48",x"d4",x"ff",x"78"),
  1623 => (x"d0",x"ff",x"78",x"71"),
  1624 => (x"78",x"e1",x"c8",x"48"),
  1625 => (x"26",x"78",x"e0",x"c0"),
  1626 => (x"5b",x"5e",x"0e",x"4f"),
  1627 => (x"4c",x"71",x"0e",x"5c"),
  1628 => (x"49",x"c3",x"f0",x"c2"),
  1629 => (x"70",x"87",x"ee",x"fa"),
  1630 => (x"aa",x"b7",x"c0",x"4a"),
  1631 => (x"87",x"e3",x"c2",x"04"),
  1632 => (x"05",x"aa",x"e0",x"c3"),
  1633 => (x"e8",x"c1",x"87",x"c9"),
  1634 => (x"78",x"c1",x"48",x"ec"),
  1635 => (x"c3",x"87",x"d4",x"c2"),
  1636 => (x"c9",x"05",x"aa",x"f0"),
  1637 => (x"e8",x"e8",x"c1",x"87"),
  1638 => (x"c1",x"78",x"c1",x"48"),
  1639 => (x"e8",x"c1",x"87",x"f5"),
  1640 => (x"c7",x"02",x"bf",x"ec"),
  1641 => (x"c2",x"4b",x"72",x"87"),
  1642 => (x"87",x"c2",x"b3",x"c0"),
  1643 => (x"9c",x"74",x"4b",x"72"),
  1644 => (x"c1",x"87",x"d1",x"05"),
  1645 => (x"1e",x"bf",x"e8",x"e8"),
  1646 => (x"bf",x"ec",x"e8",x"c1"),
  1647 => (x"fd",x"49",x"72",x"1e"),
  1648 => (x"86",x"c8",x"87",x"f8"),
  1649 => (x"bf",x"e8",x"e8",x"c1"),
  1650 => (x"87",x"e0",x"c0",x"02"),
  1651 => (x"b7",x"c4",x"49",x"73"),
  1652 => (x"ea",x"c1",x"91",x"29"),
  1653 => (x"4a",x"73",x"81",x"c8"),
  1654 => (x"92",x"c2",x"9a",x"cf"),
  1655 => (x"30",x"72",x"48",x"c1"),
  1656 => (x"ba",x"ff",x"4a",x"70"),
  1657 => (x"98",x"69",x"48",x"72"),
  1658 => (x"87",x"db",x"79",x"70"),
  1659 => (x"b7",x"c4",x"49",x"73"),
  1660 => (x"ea",x"c1",x"91",x"29"),
  1661 => (x"4a",x"73",x"81",x"c8"),
  1662 => (x"92",x"c2",x"9a",x"cf"),
  1663 => (x"30",x"72",x"48",x"c3"),
  1664 => (x"69",x"48",x"4a",x"70"),
  1665 => (x"c1",x"79",x"70",x"b0"),
  1666 => (x"c0",x"48",x"ec",x"e8"),
  1667 => (x"e8",x"e8",x"c1",x"78"),
  1668 => (x"c2",x"78",x"c0",x"48"),
  1669 => (x"f8",x"49",x"c3",x"f0"),
  1670 => (x"4a",x"70",x"87",x"cb"),
  1671 => (x"03",x"aa",x"b7",x"c0"),
  1672 => (x"c0",x"87",x"dd",x"fd"),
  1673 => (x"87",x"c8",x"fc",x"48"),
  1674 => (x"00",x"00",x"00",x"00"),
  1675 => (x"00",x"00",x"00",x"00"),
  1676 => (x"49",x"4a",x"71",x"1e"),
  1677 => (x"26",x"87",x"f2",x"fc"),
  1678 => (x"4a",x"c0",x"1e",x"4f"),
  1679 => (x"91",x"c4",x"49",x"72"),
  1680 => (x"81",x"c8",x"ea",x"c1"),
  1681 => (x"82",x"c1",x"79",x"c0"),
  1682 => (x"04",x"aa",x"b7",x"d0"),
  1683 => (x"4f",x"26",x"87",x"ee"),
  1684 => (x"5c",x"5b",x"5e",x"0e"),
  1685 => (x"4d",x"71",x"0e",x"5d"),
  1686 => (x"75",x"87",x"fa",x"f6"),
  1687 => (x"2a",x"b7",x"c4",x"4a"),
  1688 => (x"c8",x"ea",x"c1",x"92"),
  1689 => (x"cf",x"4c",x"75",x"82"),
  1690 => (x"6a",x"94",x"c2",x"9c"),
  1691 => (x"2b",x"74",x"4b",x"49"),
  1692 => (x"48",x"c2",x"9b",x"c3"),
  1693 => (x"4c",x"70",x"30",x"74"),
  1694 => (x"48",x"74",x"bc",x"ff"),
  1695 => (x"7a",x"70",x"98",x"71"),
  1696 => (x"73",x"87",x"ca",x"f6"),
  1697 => (x"87",x"e6",x"fa",x"48"),
  1698 => (x"00",x"00",x"00",x"00"),
  1699 => (x"00",x"00",x"00",x"00"),
  1700 => (x"00",x"00",x"00",x"00"),
  1701 => (x"00",x"00",x"00",x"00"),
  1702 => (x"00",x"00",x"00",x"00"),
  1703 => (x"00",x"00",x"00",x"00"),
  1704 => (x"00",x"00",x"00",x"00"),
  1705 => (x"00",x"00",x"00",x"00"),
  1706 => (x"00",x"00",x"00",x"00"),
  1707 => (x"00",x"00",x"00",x"00"),
  1708 => (x"00",x"00",x"00",x"00"),
  1709 => (x"00",x"00",x"00",x"00"),
  1710 => (x"00",x"00",x"00",x"00"),
  1711 => (x"00",x"00",x"00",x"00"),
  1712 => (x"00",x"00",x"00",x"00"),
  1713 => (x"00",x"00",x"00",x"00"),
  1714 => (x"25",x"26",x"1e",x"16"),
  1715 => (x"3e",x"3d",x"36",x"2e"),
  1716 => (x"48",x"d0",x"ff",x"1e"),
  1717 => (x"71",x"78",x"e1",x"c8"),
  1718 => (x"08",x"d4",x"ff",x"48"),
  1719 => (x"1e",x"4f",x"26",x"78"),
  1720 => (x"c8",x"48",x"d0",x"ff"),
  1721 => (x"48",x"71",x"78",x"e1"),
  1722 => (x"78",x"08",x"d4",x"ff"),
  1723 => (x"ff",x"48",x"66",x"c4"),
  1724 => (x"26",x"78",x"08",x"d4"),
  1725 => (x"4a",x"71",x"1e",x"4f"),
  1726 => (x"1e",x"49",x"66",x"c4"),
  1727 => (x"de",x"ff",x"49",x"72"),
  1728 => (x"48",x"d0",x"ff",x"87"),
  1729 => (x"26",x"78",x"e0",x"c0"),
  1730 => (x"71",x"1e",x"4f",x"26"),
  1731 => (x"1e",x"66",x"c4",x"4a"),
  1732 => (x"49",x"a2",x"e0",x"c1"),
  1733 => (x"c8",x"87",x"c8",x"ff"),
  1734 => (x"b7",x"c8",x"49",x"66"),
  1735 => (x"48",x"d4",x"ff",x"29"),
  1736 => (x"d0",x"ff",x"78",x"71"),
  1737 => (x"78",x"e0",x"c0",x"48"),
  1738 => (x"1e",x"4f",x"26",x"26"),
  1739 => (x"c3",x"4a",x"d4",x"ff"),
  1740 => (x"d0",x"ff",x"7a",x"ff"),
  1741 => (x"78",x"e1",x"c8",x"48"),
  1742 => (x"f0",x"c2",x"7a",x"de"),
  1743 => (x"49",x"7a",x"bf",x"cd"),
  1744 => (x"70",x"28",x"c8",x"48"),
  1745 => (x"d0",x"48",x"71",x"7a"),
  1746 => (x"71",x"7a",x"70",x"28"),
  1747 => (x"70",x"28",x"d8",x"48"),
  1748 => (x"48",x"d0",x"ff",x"7a"),
  1749 => (x"26",x"78",x"e0",x"c0"),
  1750 => (x"5b",x"5e",x"0e",x"4f"),
  1751 => (x"71",x"0e",x"5d",x"5c"),
  1752 => (x"cd",x"f0",x"c2",x"4c"),
  1753 => (x"74",x"4b",x"4d",x"bf"),
  1754 => (x"9b",x"66",x"d0",x"2b"),
  1755 => (x"66",x"d4",x"83",x"c1"),
  1756 => (x"87",x"c2",x"04",x"ab"),
  1757 => (x"4a",x"74",x"4b",x"c0"),
  1758 => (x"72",x"49",x"66",x"d0"),
  1759 => (x"75",x"b9",x"ff",x"31"),
  1760 => (x"72",x"48",x"73",x"99"),
  1761 => (x"48",x"4a",x"70",x"30"),
  1762 => (x"f0",x"c2",x"b0",x"71"),
  1763 => (x"da",x"fe",x"58",x"d1"),
  1764 => (x"26",x"4d",x"26",x"87"),
  1765 => (x"26",x"4b",x"26",x"4c"),
  1766 => (x"d0",x"ff",x"1e",x"4f"),
  1767 => (x"78",x"c9",x"c8",x"48"),
  1768 => (x"d4",x"ff",x"48",x"71"),
  1769 => (x"4f",x"26",x"78",x"08"),
  1770 => (x"49",x"4a",x"71",x"1e"),
  1771 => (x"d0",x"ff",x"87",x"eb"),
  1772 => (x"26",x"78",x"c8",x"48"),
  1773 => (x"1e",x"73",x"1e",x"4f"),
  1774 => (x"f0",x"c2",x"4b",x"71"),
  1775 => (x"c3",x"02",x"bf",x"dd"),
  1776 => (x"87",x"eb",x"c2",x"87"),
  1777 => (x"c8",x"48",x"d0",x"ff"),
  1778 => (x"49",x"73",x"78",x"c9"),
  1779 => (x"ff",x"b1",x"e0",x"c0"),
  1780 => (x"78",x"71",x"48",x"d4"),
  1781 => (x"48",x"d1",x"f0",x"c2"),
  1782 => (x"66",x"c8",x"78",x"c0"),
  1783 => (x"c3",x"87",x"c5",x"02"),
  1784 => (x"87",x"c2",x"49",x"ff"),
  1785 => (x"f0",x"c2",x"49",x"c0"),
  1786 => (x"66",x"cc",x"59",x"d9"),
  1787 => (x"c5",x"87",x"c6",x"02"),
  1788 => (x"c4",x"4a",x"d5",x"d5"),
  1789 => (x"ff",x"ff",x"cf",x"87"),
  1790 => (x"dd",x"f0",x"c2",x"4a"),
  1791 => (x"dd",x"f0",x"c2",x"5a"),
  1792 => (x"c4",x"78",x"c1",x"48"),
  1793 => (x"26",x"4d",x"26",x"87"),
  1794 => (x"26",x"4b",x"26",x"4c"),
  1795 => (x"5b",x"5e",x"0e",x"4f"),
  1796 => (x"71",x"0e",x"5d",x"5c"),
  1797 => (x"d9",x"f0",x"c2",x"4a"),
  1798 => (x"9a",x"72",x"4c",x"bf"),
  1799 => (x"49",x"87",x"cb",x"02"),
  1800 => (x"ee",x"c1",x"91",x"c8"),
  1801 => (x"83",x"71",x"4b",x"eb"),
  1802 => (x"f2",x"c1",x"87",x"c4"),
  1803 => (x"4d",x"c0",x"4b",x"eb"),
  1804 => (x"99",x"74",x"49",x"13"),
  1805 => (x"bf",x"d5",x"f0",x"c2"),
  1806 => (x"48",x"d4",x"ff",x"b9"),
  1807 => (x"b7",x"c1",x"78",x"71"),
  1808 => (x"b7",x"c8",x"85",x"2c"),
  1809 => (x"87",x"e8",x"04",x"ad"),
  1810 => (x"bf",x"d1",x"f0",x"c2"),
  1811 => (x"c2",x"80",x"c8",x"48"),
  1812 => (x"fe",x"58",x"d5",x"f0"),
  1813 => (x"73",x"1e",x"87",x"ef"),
  1814 => (x"13",x"4b",x"71",x"1e"),
  1815 => (x"cb",x"02",x"9a",x"4a"),
  1816 => (x"fe",x"49",x"72",x"87"),
  1817 => (x"4a",x"13",x"87",x"e7"),
  1818 => (x"87",x"f5",x"05",x"9a"),
  1819 => (x"1e",x"87",x"da",x"fe"),
  1820 => (x"bf",x"d1",x"f0",x"c2"),
  1821 => (x"d1",x"f0",x"c2",x"49"),
  1822 => (x"78",x"a1",x"c1",x"48"),
  1823 => (x"a9",x"b7",x"c0",x"c4"),
  1824 => (x"ff",x"87",x"db",x"03"),
  1825 => (x"f0",x"c2",x"48",x"d4"),
  1826 => (x"c2",x"78",x"bf",x"d5"),
  1827 => (x"49",x"bf",x"d1",x"f0"),
  1828 => (x"48",x"d1",x"f0",x"c2"),
  1829 => (x"c4",x"78",x"a1",x"c1"),
  1830 => (x"04",x"a9",x"b7",x"c0"),
  1831 => (x"d0",x"ff",x"87",x"e5"),
  1832 => (x"c2",x"78",x"c8",x"48"),
  1833 => (x"c0",x"48",x"dd",x"f0"),
  1834 => (x"00",x"4f",x"26",x"78"),
  1835 => (x"00",x"00",x"00",x"00"),
  1836 => (x"00",x"00",x"00",x"00"),
  1837 => (x"5f",x"5f",x"00",x"00"),
  1838 => (x"00",x"00",x"00",x"00"),
  1839 => (x"03",x"00",x"03",x"03"),
  1840 => (x"14",x"00",x"00",x"03"),
  1841 => (x"7f",x"14",x"7f",x"7f"),
  1842 => (x"00",x"00",x"14",x"7f"),
  1843 => (x"6b",x"6b",x"2e",x"24"),
  1844 => (x"4c",x"00",x"12",x"3a"),
  1845 => (x"6c",x"18",x"36",x"6a"),
  1846 => (x"30",x"00",x"32",x"56"),
  1847 => (x"77",x"59",x"4f",x"7e"),
  1848 => (x"00",x"40",x"68",x"3a"),
  1849 => (x"03",x"07",x"04",x"00"),
  1850 => (x"00",x"00",x"00",x"00"),
  1851 => (x"63",x"3e",x"1c",x"00"),
  1852 => (x"00",x"00",x"00",x"41"),
  1853 => (x"3e",x"63",x"41",x"00"),
  1854 => (x"08",x"00",x"00",x"1c"),
  1855 => (x"1c",x"1c",x"3e",x"2a"),
  1856 => (x"00",x"08",x"2a",x"3e"),
  1857 => (x"3e",x"3e",x"08",x"08"),
  1858 => (x"00",x"00",x"08",x"08"),
  1859 => (x"60",x"e0",x"80",x"00"),
  1860 => (x"00",x"00",x"00",x"00"),
  1861 => (x"08",x"08",x"08",x"08"),
  1862 => (x"00",x"00",x"08",x"08"),
  1863 => (x"60",x"60",x"00",x"00"),
  1864 => (x"40",x"00",x"00",x"00"),
  1865 => (x"0c",x"18",x"30",x"60"),
  1866 => (x"00",x"01",x"03",x"06"),
  1867 => (x"4d",x"59",x"7f",x"3e"),
  1868 => (x"00",x"00",x"3e",x"7f"),
  1869 => (x"7f",x"7f",x"06",x"04"),
  1870 => (x"00",x"00",x"00",x"00"),
  1871 => (x"59",x"71",x"63",x"42"),
  1872 => (x"00",x"00",x"46",x"4f"),
  1873 => (x"49",x"49",x"63",x"22"),
  1874 => (x"18",x"00",x"36",x"7f"),
  1875 => (x"7f",x"13",x"16",x"1c"),
  1876 => (x"00",x"00",x"10",x"7f"),
  1877 => (x"45",x"45",x"67",x"27"),
  1878 => (x"00",x"00",x"39",x"7d"),
  1879 => (x"49",x"4b",x"7e",x"3c"),
  1880 => (x"00",x"00",x"30",x"79"),
  1881 => (x"79",x"71",x"01",x"01"),
  1882 => (x"00",x"00",x"07",x"0f"),
  1883 => (x"49",x"49",x"7f",x"36"),
  1884 => (x"00",x"00",x"36",x"7f"),
  1885 => (x"69",x"49",x"4f",x"06"),
  1886 => (x"00",x"00",x"1e",x"3f"),
  1887 => (x"66",x"66",x"00",x"00"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"66",x"e6",x"80",x"00"),
  1890 => (x"00",x"00",x"00",x"00"),
  1891 => (x"14",x"14",x"08",x"08"),
  1892 => (x"00",x"00",x"22",x"22"),
  1893 => (x"14",x"14",x"14",x"14"),
  1894 => (x"00",x"00",x"14",x"14"),
  1895 => (x"14",x"14",x"22",x"22"),
  1896 => (x"00",x"00",x"08",x"08"),
  1897 => (x"59",x"51",x"03",x"02"),
  1898 => (x"3e",x"00",x"06",x"0f"),
  1899 => (x"55",x"5d",x"41",x"7f"),
  1900 => (x"00",x"00",x"1e",x"1f"),
  1901 => (x"09",x"09",x"7f",x"7e"),
  1902 => (x"00",x"00",x"7e",x"7f"),
  1903 => (x"49",x"49",x"7f",x"7f"),
  1904 => (x"00",x"00",x"36",x"7f"),
  1905 => (x"41",x"63",x"3e",x"1c"),
  1906 => (x"00",x"00",x"41",x"41"),
  1907 => (x"63",x"41",x"7f",x"7f"),
  1908 => (x"00",x"00",x"1c",x"3e"),
  1909 => (x"49",x"49",x"7f",x"7f"),
  1910 => (x"00",x"00",x"41",x"41"),
  1911 => (x"09",x"09",x"7f",x"7f"),
  1912 => (x"00",x"00",x"01",x"01"),
  1913 => (x"49",x"41",x"7f",x"3e"),
  1914 => (x"00",x"00",x"7a",x"7b"),
  1915 => (x"08",x"08",x"7f",x"7f"),
  1916 => (x"00",x"00",x"7f",x"7f"),
  1917 => (x"7f",x"7f",x"41",x"00"),
  1918 => (x"00",x"00",x"00",x"41"),
  1919 => (x"40",x"40",x"60",x"20"),
  1920 => (x"7f",x"00",x"3f",x"7f"),
  1921 => (x"36",x"1c",x"08",x"7f"),
  1922 => (x"00",x"00",x"41",x"63"),
  1923 => (x"40",x"40",x"7f",x"7f"),
  1924 => (x"7f",x"00",x"40",x"40"),
  1925 => (x"06",x"0c",x"06",x"7f"),
  1926 => (x"7f",x"00",x"7f",x"7f"),
  1927 => (x"18",x"0c",x"06",x"7f"),
  1928 => (x"00",x"00",x"7f",x"7f"),
  1929 => (x"41",x"41",x"7f",x"3e"),
  1930 => (x"00",x"00",x"3e",x"7f"),
  1931 => (x"09",x"09",x"7f",x"7f"),
  1932 => (x"3e",x"00",x"06",x"0f"),
  1933 => (x"7f",x"61",x"41",x"7f"),
  1934 => (x"00",x"00",x"40",x"7e"),
  1935 => (x"19",x"09",x"7f",x"7f"),
  1936 => (x"00",x"00",x"66",x"7f"),
  1937 => (x"59",x"4d",x"6f",x"26"),
  1938 => (x"00",x"00",x"32",x"7b"),
  1939 => (x"7f",x"7f",x"01",x"01"),
  1940 => (x"00",x"00",x"01",x"01"),
  1941 => (x"40",x"40",x"7f",x"3f"),
  1942 => (x"00",x"00",x"3f",x"7f"),
  1943 => (x"70",x"70",x"3f",x"0f"),
  1944 => (x"7f",x"00",x"0f",x"3f"),
  1945 => (x"30",x"18",x"30",x"7f"),
  1946 => (x"41",x"00",x"7f",x"7f"),
  1947 => (x"1c",x"1c",x"36",x"63"),
  1948 => (x"01",x"41",x"63",x"36"),
  1949 => (x"7c",x"7c",x"06",x"03"),
  1950 => (x"61",x"01",x"03",x"06"),
  1951 => (x"47",x"4d",x"59",x"71"),
  1952 => (x"00",x"00",x"41",x"43"),
  1953 => (x"41",x"7f",x"7f",x"00"),
  1954 => (x"01",x"00",x"00",x"41"),
  1955 => (x"18",x"0c",x"06",x"03"),
  1956 => (x"00",x"40",x"60",x"30"),
  1957 => (x"7f",x"41",x"41",x"00"),
  1958 => (x"08",x"00",x"00",x"7f"),
  1959 => (x"06",x"03",x"06",x"0c"),
  1960 => (x"80",x"00",x"08",x"0c"),
  1961 => (x"80",x"80",x"80",x"80"),
  1962 => (x"00",x"00",x"80",x"80"),
  1963 => (x"07",x"03",x"00",x"00"),
  1964 => (x"00",x"00",x"00",x"04"),
  1965 => (x"54",x"54",x"74",x"20"),
  1966 => (x"00",x"00",x"78",x"7c"),
  1967 => (x"44",x"44",x"7f",x"7f"),
  1968 => (x"00",x"00",x"38",x"7c"),
  1969 => (x"44",x"44",x"7c",x"38"),
  1970 => (x"00",x"00",x"00",x"44"),
  1971 => (x"44",x"44",x"7c",x"38"),
  1972 => (x"00",x"00",x"7f",x"7f"),
  1973 => (x"54",x"54",x"7c",x"38"),
  1974 => (x"00",x"00",x"18",x"5c"),
  1975 => (x"05",x"7f",x"7e",x"04"),
  1976 => (x"00",x"00",x"00",x"05"),
  1977 => (x"a4",x"a4",x"bc",x"18"),
  1978 => (x"00",x"00",x"7c",x"fc"),
  1979 => (x"04",x"04",x"7f",x"7f"),
  1980 => (x"00",x"00",x"78",x"7c"),
  1981 => (x"7d",x"3d",x"00",x"00"),
  1982 => (x"00",x"00",x"00",x"40"),
  1983 => (x"fd",x"80",x"80",x"80"),
  1984 => (x"00",x"00",x"00",x"7d"),
  1985 => (x"38",x"10",x"7f",x"7f"),
  1986 => (x"00",x"00",x"44",x"6c"),
  1987 => (x"7f",x"3f",x"00",x"00"),
  1988 => (x"7c",x"00",x"00",x"40"),
  1989 => (x"0c",x"18",x"0c",x"7c"),
  1990 => (x"00",x"00",x"78",x"7c"),
  1991 => (x"04",x"04",x"7c",x"7c"),
  1992 => (x"00",x"00",x"78",x"7c"),
  1993 => (x"44",x"44",x"7c",x"38"),
  1994 => (x"00",x"00",x"38",x"7c"),
  1995 => (x"24",x"24",x"fc",x"fc"),
  1996 => (x"00",x"00",x"18",x"3c"),
  1997 => (x"24",x"24",x"3c",x"18"),
  1998 => (x"00",x"00",x"fc",x"fc"),
  1999 => (x"04",x"04",x"7c",x"7c"),
  2000 => (x"00",x"00",x"08",x"0c"),
  2001 => (x"54",x"54",x"5c",x"48"),
  2002 => (x"00",x"00",x"20",x"74"),
  2003 => (x"44",x"7f",x"3f",x"04"),
  2004 => (x"00",x"00",x"00",x"44"),
  2005 => (x"40",x"40",x"7c",x"3c"),
  2006 => (x"00",x"00",x"7c",x"7c"),
  2007 => (x"60",x"60",x"3c",x"1c"),
  2008 => (x"3c",x"00",x"1c",x"3c"),
  2009 => (x"60",x"30",x"60",x"7c"),
  2010 => (x"44",x"00",x"3c",x"7c"),
  2011 => (x"38",x"10",x"38",x"6c"),
  2012 => (x"00",x"00",x"44",x"6c"),
  2013 => (x"60",x"e0",x"bc",x"1c"),
  2014 => (x"00",x"00",x"1c",x"3c"),
  2015 => (x"5c",x"74",x"64",x"44"),
  2016 => (x"00",x"00",x"44",x"4c"),
  2017 => (x"77",x"3e",x"08",x"08"),
  2018 => (x"00",x"00",x"41",x"41"),
  2019 => (x"7f",x"7f",x"00",x"00"),
  2020 => (x"00",x"00",x"00",x"00"),
  2021 => (x"3e",x"77",x"41",x"41"),
  2022 => (x"02",x"00",x"08",x"08"),
  2023 => (x"02",x"03",x"01",x"01"),
  2024 => (x"7f",x"00",x"01",x"02"),
  2025 => (x"7f",x"7f",x"7f",x"7f"),
  2026 => (x"08",x"00",x"7f",x"7f"),
  2027 => (x"3e",x"1c",x"1c",x"08"),
  2028 => (x"7f",x"7f",x"7f",x"3e"),
  2029 => (x"1c",x"3e",x"3e",x"7f"),
  2030 => (x"00",x"08",x"08",x"1c"),
  2031 => (x"7c",x"7c",x"18",x"10"),
  2032 => (x"00",x"00",x"10",x"18"),
  2033 => (x"7c",x"7c",x"30",x"10"),
  2034 => (x"10",x"00",x"10",x"30"),
  2035 => (x"78",x"60",x"60",x"30"),
  2036 => (x"42",x"00",x"06",x"1e"),
  2037 => (x"3c",x"18",x"3c",x"66"),
  2038 => (x"78",x"00",x"42",x"66"),
  2039 => (x"c6",x"c2",x"6a",x"38"),
  2040 => (x"60",x"00",x"38",x"6c"),
  2041 => (x"00",x"60",x"00",x"00"),
  2042 => (x"0e",x"00",x"60",x"00"),
  2043 => (x"5d",x"5c",x"5b",x"5e"),
  2044 => (x"4c",x"71",x"1e",x"0e"),
  2045 => (x"bf",x"ee",x"f0",x"c2"),
  2046 => (x"c0",x"4b",x"c0",x"4d"),
  2047 => (x"02",x"ab",x"74",x"1e"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

